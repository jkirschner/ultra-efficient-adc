magic
tech scmos
timestamp 1355432294
<< ntransistor >>
rect 17 -7 20 3
<< ptransistor >>
rect 17 15 20 35
<< ndiffusion >>
rect 14 -3 17 3
rect 16 -7 17 -3
rect 20 -1 21 3
rect 20 -7 23 -1
<< pdiffusion >>
rect 14 34 17 35
rect 15 24 17 34
rect 14 15 17 24
rect 20 20 23 35
rect 20 16 21 20
rect 20 15 23 16
<< ndcontact >>
rect 12 -7 16 -3
rect 21 -1 25 3
<< pdcontact >>
rect 11 24 15 34
rect 21 16 25 20
<< psubstratepcontact >>
rect 26 -18 30 -14
<< nsubstratencontact >>
rect 31 33 35 37
<< polysilicon >>
rect 17 35 20 37
rect 17 10 20 15
rect 18 6 20 10
rect 17 3 20 6
rect 17 -9 20 -7
<< polycontact >>
rect 14 6 18 10
<< metal1 >>
rect -5 37 43 41
rect -5 34 31 37
rect -5 24 11 34
rect 15 33 31 34
rect 35 33 43 37
rect 15 24 43 33
rect -5 23 43 24
rect 21 10 25 16
rect -5 6 14 10
rect 21 6 43 10
rect 21 3 25 6
rect -5 -7 12 -4
rect 16 -7 43 -4
rect -5 -14 43 -7
rect -5 -18 26 -14
rect 30 -18 43 -14
rect -5 -23 43 -18
<< labels >>
rlabel metal1 -4 8 -4 8 3 In
rlabel metal1 42 8 42 8 7 Out
rlabel metal1 4 -21 4 -21 1 Gnd
rlabel metal1 4 35 4 35 1 Vdd
<< end >>
