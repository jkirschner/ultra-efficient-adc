* SPICE3 file created from PulseWidthControl_Layout.ext - technology: scmos

M1000 a_3_28# a_1_26# Vpos Vpos pfet w=1.8u l=0.6u
+ ad=4.68p pd=13.2u as=30.06p ps=61.2u 
M1001 a_19_77# OutB a_18_41# Vpos pfet w=1.8u l=0.6u
+ ad=2.34p pd=6.6u as=5.4p ps=13.8u 
M1002 a_1_26# Din Vpos Vpos pfet w=1.8u l=0.6u
+ ad=2.34p pd=6.6u as=0p ps=0u 
M1003 Vneg Out Din Vneg nfet w=4.5u l=2.4u
+ ad=27.09p pd=61.2u as=6.75p ps=12u 
M1004 a_1_26# Din Vneg Vneg nfet w=0.9u l=0.6u
+ ad=1.71p pd=5.4u as=0p ps=0u 
M1005 Vpos a_30_70# a_32_67# Vpos pfet w=7.2u l=3.6u
+ ad=0p pd=0u as=10.62p ps=22.8u 
M1006 Vpos Vpw2 a_61_55# Vpos pfet w=4.8u l=1.8u
+ ad=0p pd=0u as=12.24p ps=25.8u 
M1007 Vpos Reset a_87_54# Vpos pfet w=1.8u l=0.6u
+ ad=0p pd=0u as=5.58p ps=13.8u 
M1008 OutB Out Vpos Vpos pfet w=3.6u l=0.6u
+ ad=3.96p pd=10.2u as=0p ps=0u 
M1009 a_18_41# Out a_3_28# Vpos pfet w=1.8u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1010 a_32_67# a_32_52# a_18_41# Vpos pfet w=1.2u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1011 a_18_41# OutB a_3_28# Vneg nfet w=0.9u l=0.6u
+ ad=3.42p pd=10.8u as=3.42p ps=10.8u 
M1012 Vpos a_18_41# a_32_52# Vpos pfet w=1.8u l=0.6u
+ ad=0p pd=0u as=2.34p ps=6.6u 
M1013 a_30_70# a_32_52# a_61_55# Vpos pfet w=1.8u l=0.9u
+ ad=3.24p pd=7.2u as=0p ps=0u 
M1014 a_61_55# a_32_52# a_30_70# Vpos pfet w=1.8u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1015 a_19_77# Out a_18_41# Vneg nfet w=0.9u l=0.6u
+ ad=9.18p pd=15u as=0p ps=0u 
M1016 a_3_28# a_1_26# Vneg Vneg nfet w=0.9u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1017 Vneg Vpw1 a_19_77# Vneg nfet w=4.5u l=2.4u
+ ad=0p pd=0u as=0p ps=0u 
M1018 a_32_52# a_18_41# Vneg Vneg nfet w=0.9u l=0.6u
+ ad=1.71p pd=5.4u as=0p ps=0u 
M1019 a_30_70# a_32_52# Vneg Vneg nfet w=0.9u l=0.9u
+ ad=1.98p pd=6u as=0p ps=0u 
M1020 Vneg a_32_52# a_30_70# Vneg nfet w=0.9u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1021 Out a_32_52# a_87_54# Vpos pfet w=1.8u l=0.6u
+ ad=2.34p pd=6.6u as=0p ps=0u 
M1022 Out a_32_52# a_78_28# Vneg nfet w=0.9u l=0.6u
+ ad=3.69p pd=8.4u as=3.78p ps=11.4u 
M1023 OutB Out Vneg Vneg nfet w=1.8u l=0.6u
+ ad=2.7p pd=7.2u as=0p ps=0u 
M1024 Out Reset Vneg Vneg nfet w=0.9u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1025 a_78_28# ResetB Vneg Vneg nfet w=0.9u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
