magic
tech scmos
timestamp 1355369771
<< nwell >>
rect -27 53 122 93
rect 13 51 122 53
rect 29 50 122 51
rect 39 49 122 50
rect 78 48 122 49
<< pwell >>
rect -27 51 13 53
rect -27 50 29 51
rect -27 49 39 50
rect -27 48 78 49
rect -27 20 122 48
<< ntransistor >>
rect -15 29 -7 44
rect 0 44 2 47
rect 16 41 18 44
rect 24 34 26 37
rect 1 28 3 31
rect 36 28 44 43
rect 50 38 52 41
rect 66 38 69 41
rect 75 38 78 41
rect 92 38 94 41
rect 106 34 112 36
rect 95 31 98 33
rect 76 28 78 31
<< ptransistor >>
rect 4 73 6 79
rect 19 75 25 77
rect 0 60 2 66
rect 32 70 56 82
rect 67 76 83 82
rect 93 71 95 77
rect 102 69 104 81
rect 24 57 26 63
rect 32 57 35 61
rect 49 55 51 61
rect 66 55 69 61
rect 75 55 78 61
rect 92 54 94 60
<< ndiffusion >>
rect -16 29 -15 44
rect -7 41 -6 44
rect -2 44 0 47
rect 2 44 3 47
rect -2 41 -1 44
rect -7 39 -1 41
rect 15 41 16 44
rect 18 41 19 44
rect -7 31 -3 39
rect 33 37 36 43
rect 23 34 24 37
rect 26 34 27 37
rect -7 29 -6 31
rect 0 28 1 31
rect 3 28 4 31
rect 35 28 36 37
rect 44 41 49 43
rect 44 30 45 41
rect 49 38 50 41
rect 52 38 53 41
rect 65 38 66 41
rect 69 38 70 41
rect 74 38 75 41
rect 78 38 79 41
rect 91 38 92 41
rect 94 38 95 41
rect 106 41 110 42
rect 110 37 112 39
rect 106 36 112 37
rect 95 33 98 34
rect 106 33 112 34
rect 44 28 49 30
rect 75 28 76 31
rect 78 28 79 31
rect 95 30 98 31
rect 99 26 100 30
rect 110 31 112 33
<< pdiffusion >>
rect 32 83 33 85
rect 55 83 56 85
rect 32 82 56 83
rect 81 83 83 87
rect 67 82 83 83
rect 1 77 4 79
rect 3 73 4 77
rect 6 77 9 79
rect 19 78 21 80
rect 19 77 25 78
rect 6 73 7 77
rect -3 64 0 66
rect -1 60 0 64
rect 2 64 5 66
rect 2 60 3 64
rect 19 74 25 75
rect 23 72 25 74
rect 99 77 102 81
rect 67 75 83 76
rect 89 75 93 77
rect 67 73 68 75
rect 32 69 56 70
rect 82 73 83 75
rect 91 71 93 75
rect 95 73 96 77
rect 100 73 102 77
rect 95 71 102 73
rect 32 67 38 69
rect 36 65 38 67
rect 49 67 56 69
rect 99 69 102 71
rect 104 77 107 81
rect 104 73 105 77
rect 104 69 107 73
rect 21 61 24 63
rect 23 57 24 61
rect 26 59 27 63
rect 31 59 32 61
rect 26 57 32 59
rect 35 57 36 61
rect 48 57 49 61
rect 46 55 49 57
rect 51 57 52 61
rect 51 55 54 57
rect 65 55 66 61
rect 69 59 75 61
rect 69 55 70 59
rect 74 55 75 59
rect 78 55 79 61
rect 91 54 92 60
rect 94 58 97 60
rect 94 54 95 58
<< ndcontact >>
rect -20 29 -16 44
rect -6 41 -2 47
rect 3 43 7 47
rect 11 40 15 44
rect 19 41 23 45
rect 19 33 23 37
rect -6 27 0 31
rect 4 27 8 31
rect 27 28 35 37
rect 45 30 49 41
rect 53 37 57 41
rect 61 35 65 41
rect 70 37 74 41
rect 79 38 83 42
rect 87 36 91 41
rect 95 34 100 41
rect 106 37 110 41
rect 71 27 75 31
rect 79 27 83 31
rect 95 26 99 30
rect 106 29 110 33
<< pdcontact >>
rect 33 83 55 87
rect 67 83 81 87
rect -1 73 3 77
rect 21 78 25 82
rect 7 73 11 77
rect -5 60 -1 64
rect 3 60 7 64
rect 19 70 23 74
rect 68 71 82 75
rect 87 71 91 75
rect 96 73 100 77
rect 38 65 49 69
rect 105 73 109 77
rect 19 57 23 61
rect 27 59 31 63
rect 36 57 40 61
rect 44 57 48 61
rect 52 57 56 61
rect 61 55 65 61
rect 70 55 74 59
rect 79 55 83 61
rect 87 54 91 60
rect 95 54 99 58
<< psubstratepdiff >>
rect 61 27 65 31
<< nsubstratendiff >>
rect -5 73 -1 77
<< psubstratepcontact >>
rect 57 27 61 31
<< nsubstratencontact >>
rect -9 73 -5 77
<< polysilicon >>
rect 4 79 6 81
rect 15 77 18 81
rect 13 75 19 77
rect 25 75 27 77
rect 4 71 6 73
rect 0 66 2 68
rect 0 47 2 60
rect -15 44 -7 46
rect 0 42 2 44
rect 13 46 18 75
rect 30 70 32 82
rect 56 73 58 82
rect 65 76 67 82
rect 83 78 84 82
rect 102 81 104 83
rect 83 76 85 78
rect 93 77 95 79
rect 56 70 57 73
rect 93 68 95 71
rect 84 66 95 68
rect 102 68 104 69
rect 102 66 103 68
rect 24 63 26 65
rect 32 61 35 63
rect 49 61 51 63
rect 66 61 69 63
rect 75 61 78 63
rect 16 44 18 46
rect 24 56 26 57
rect 24 44 27 56
rect 32 55 35 57
rect 32 54 44 55
rect 32 52 40 54
rect 49 53 51 55
rect 49 48 52 53
rect 66 51 69 55
rect 75 51 78 55
rect 65 50 78 51
rect 16 39 18 41
rect 24 37 26 44
rect 36 43 44 45
rect 66 46 76 50
rect 1 31 3 34
rect -15 27 -7 29
rect 1 26 3 28
rect 24 29 26 34
rect 22 25 26 29
rect 50 41 52 44
rect 66 45 78 46
rect 66 41 69 45
rect 75 41 78 45
rect 50 36 52 38
rect 66 36 69 38
rect 75 36 78 38
rect 84 35 86 66
rect 92 60 94 62
rect 92 50 94 54
rect 92 41 94 46
rect 102 43 105 47
rect 92 36 94 38
rect 84 33 89 35
rect 103 36 105 43
rect 103 34 106 36
rect 112 34 114 36
rect 76 31 78 33
rect 84 31 95 33
rect 98 31 100 33
rect 36 26 44 28
rect 76 24 78 28
rect 84 29 94 31
rect 88 24 94 29
rect 92 23 94 24
<< polycontact >>
rect 3 81 7 85
rect 14 81 18 85
rect -4 51 0 55
rect 84 78 88 82
rect 57 69 61 73
rect 40 50 44 54
rect 1 34 5 38
rect 26 40 30 44
rect 48 44 52 48
rect 62 46 66 50
rect 76 46 80 50
rect -13 23 -9 27
rect 103 64 107 68
rect 90 46 94 50
rect 98 43 102 47
rect 22 21 26 25
rect 38 22 42 26
rect 75 20 79 24
rect 88 20 92 24
<< metal1 >>
rect -27 77 -1 89
rect 55 83 67 87
rect 25 78 29 82
rect 84 82 88 93
rect 96 84 122 89
rect 96 82 102 84
rect 100 78 102 82
rect 23 77 29 78
rect -27 73 -9 77
rect -5 68 -1 77
rect 11 73 14 74
rect 7 71 14 73
rect -27 51 -4 55
rect -27 47 -16 51
rect 3 47 7 60
rect 10 61 14 71
rect 26 70 29 77
rect 96 77 102 78
rect 19 67 23 70
rect 100 73 102 77
rect 112 73 122 84
rect 19 64 31 67
rect 27 63 31 64
rect 10 57 19 61
rect 73 65 77 71
rect 38 61 41 65
rect 10 56 15 57
rect -20 44 -16 47
rect -6 35 -3 41
rect 1 40 7 43
rect 11 44 15 56
rect 28 54 31 59
rect 40 57 41 61
rect 61 62 82 65
rect 61 61 65 62
rect 45 54 48 57
rect 79 61 82 62
rect 87 60 90 71
rect 1 38 5 40
rect 11 31 15 40
rect 19 51 37 54
rect 19 45 22 51
rect 19 37 23 41
rect 34 47 37 51
rect 44 51 58 54
rect 70 51 73 55
rect 103 58 106 64
rect 99 57 106 58
rect 99 54 122 57
rect 55 50 58 51
rect 34 44 48 47
rect 55 46 62 50
rect 97 52 122 54
rect 55 41 58 46
rect 70 41 73 47
rect 80 46 90 50
rect 97 47 101 52
rect 97 43 98 47
rect 106 45 122 46
rect 97 42 101 43
rect 8 27 15 31
rect 35 34 39 37
rect 57 37 58 41
rect 95 41 101 42
rect 110 41 122 45
rect 61 34 65 35
rect 49 30 51 34
rect 45 27 51 30
rect 55 31 68 34
rect 87 31 91 36
rect 55 27 57 31
rect 61 27 71 31
rect 83 27 91 31
rect 97 30 106 31
rect 103 29 106 30
rect 103 26 110 29
rect -9 23 22 24
rect -13 21 22 23
rect 38 20 42 22
<< m2contact >>
rect 14 85 18 89
rect 7 81 11 85
rect 43 79 47 83
rect 96 78 100 82
rect -5 64 -1 68
rect 3 64 7 68
rect 29 70 33 74
rect 61 69 65 73
rect 105 77 109 81
rect 52 61 56 65
rect -6 31 -2 35
rect 26 44 30 48
rect 95 58 99 62
rect 69 47 73 51
rect 35 37 39 41
rect 106 41 110 45
rect 79 34 83 38
rect 51 27 55 34
rect 99 26 103 30
<< metal2 >>
rect 18 86 109 89
rect 3 68 7 85
rect 21 82 43 83
rect 14 79 43 82
rect 47 82 100 83
rect 47 79 96 82
rect 14 78 96 79
rect 105 81 109 86
rect 10 77 96 78
rect 10 74 26 77
rect 36 76 96 77
rect -5 61 -1 64
rect 10 61 18 74
rect -5 57 18 61
rect -5 56 17 57
rect 29 54 33 70
rect 43 67 53 76
rect 105 73 109 77
rect 43 65 56 67
rect 43 61 52 65
rect 43 57 56 61
rect 61 59 65 69
rect 61 55 73 59
rect 20 51 33 54
rect 69 51 73 55
rect 20 40 23 51
rect 30 45 66 48
rect 63 44 66 45
rect 95 44 99 58
rect 105 45 110 73
rect 63 41 99 44
rect 31 40 35 41
rect -27 35 -22 39
rect 20 37 35 40
rect -27 31 -6 35
rect -2 31 51 34
rect -27 27 51 31
rect 55 33 83 34
rect 112 33 122 38
rect 55 30 122 33
rect 55 27 99 30
rect 95 26 99 27
rect 103 26 122 30
<< labels >>
rlabel metal1 84 92 88 93 5 Vpw2
rlabel metal1 99 50 99 50 1 Out
rlabel metal2 108 50 108 50 7 OutB
rlabel ndcontact 47 30 47 30 7 Vneg
rlabel metal1 -11 22 -11 22 1 Out
rlabel polysilicon 25 30 25 30 1 Out
rlabel metal1 121 41 122 46 7 OutB
rlabel metal1 121 52 122 57 7 Out
rlabel metal2 121 26 122 38 7 Vneg
rlabel metal1 121 73 122 89 7 Vpos
rlabel metal1 -27 73 -26 89 3 Vpos
rlabel metal2 -27 27 -26 39 3 Vneg
rlabel metal1 -27 47 -26 55 3 Din
rlabel metal1 38 20 42 21 1 Vpw1
rlabel polycontact 88 20 92 21 1 Reset
rlabel polycontact 75 20 79 21 1 ResetB
<< end >>
