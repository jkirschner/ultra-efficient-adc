magic
tech scmos
timestamp 1355437586
<< ntransistor >>
rect -18 -49 -5 -42
rect 1 -49 14 -42
rect 20 -47 47 -44
rect 60 -48 73 -21
rect 117 -48 130 -21
rect 143 -47 170 -44
rect 176 -49 189 -42
rect 195 -49 208 -42
rect 60 -59 73 -52
rect 79 -59 92 -52
rect 98 -59 111 -52
rect 117 -59 130 -52
<< ptransistor >>
rect 25 29 38 56
rect 44 29 57 56
rect 133 29 146 56
rect 152 29 165 56
rect 6 -9 19 18
rect 25 -9 38 18
rect 44 -9 47 18
rect 60 3 73 9
rect 79 -9 92 18
rect 98 -9 111 18
rect 117 3 130 9
rect 143 -9 146 18
rect 152 -9 165 18
rect 171 -9 184 18
<< ndiffusion >>
rect 57 -22 60 -21
rect 59 -26 60 -22
rect -21 -44 -18 -42
rect -19 -48 -18 -44
rect -21 -49 -18 -48
rect -5 -46 -4 -42
rect 0 -46 1 -42
rect -5 -49 1 -46
rect 14 -44 17 -42
rect 14 -48 15 -44
rect 19 -47 20 -44
rect 47 -47 48 -44
rect 14 -49 17 -48
rect 57 -48 60 -26
rect 73 -42 76 -21
rect 114 -42 117 -21
rect 73 -46 74 -42
rect 116 -46 117 -42
rect 73 -48 76 -46
rect 114 -48 117 -46
rect 130 -22 133 -21
rect 130 -26 131 -22
rect 130 -48 133 -26
rect 173 -44 176 -42
rect 142 -47 143 -44
rect 170 -47 171 -44
rect 175 -48 176 -44
rect 173 -49 176 -48
rect 189 -46 190 -42
rect 194 -46 195 -42
rect 189 -49 195 -46
rect 208 -44 211 -42
rect 208 -48 209 -44
rect 208 -49 211 -48
rect 57 -54 60 -52
rect 59 -58 60 -54
rect 57 -59 60 -58
rect 73 -53 79 -52
rect 73 -57 74 -53
rect 78 -57 79 -53
rect 73 -59 79 -57
rect 92 -56 93 -52
rect 97 -56 98 -52
rect 92 -59 98 -56
rect 111 -53 117 -52
rect 111 -57 112 -53
rect 116 -57 117 -53
rect 111 -59 117 -57
rect 130 -54 133 -52
rect 130 -58 131 -54
rect 130 -59 133 -58
<< pdiffusion >>
rect 22 55 25 56
rect 24 47 25 55
rect 22 29 25 47
rect 38 34 44 56
rect 38 30 39 34
rect 43 30 44 34
rect 38 29 44 30
rect 57 55 60 56
rect 130 55 133 56
rect 57 47 58 55
rect 132 47 133 55
rect 57 29 60 47
rect 130 29 133 47
rect 146 34 152 56
rect 146 30 147 34
rect 151 30 152 34
rect 146 29 152 30
rect 165 54 168 56
rect 165 47 166 54
rect 165 29 168 47
rect 3 17 6 18
rect 5 13 6 17
rect 3 -9 6 13
rect 19 17 25 18
rect 19 -7 20 17
rect 24 -7 25 17
rect 19 -9 25 -7
rect 38 17 44 18
rect 38 13 39 17
rect 43 13 44 17
rect 38 -9 44 13
rect 47 17 50 18
rect 47 13 48 17
rect 47 -9 50 13
rect 76 9 79 18
rect 57 7 60 9
rect 59 3 60 7
rect 73 5 74 9
rect 78 5 79 9
rect 73 3 79 5
rect 76 -9 79 3
rect 92 -3 98 18
rect 92 -7 93 -3
rect 97 -7 98 -3
rect 92 -9 98 -7
rect 111 9 114 18
rect 140 17 143 18
rect 142 13 143 17
rect 111 5 112 9
rect 116 5 117 9
rect 111 3 117 5
rect 130 7 133 9
rect 130 3 131 7
rect 111 -9 114 3
rect 140 -9 143 13
rect 146 17 152 18
rect 146 13 147 17
rect 151 13 152 17
rect 146 -9 152 13
rect 165 17 171 18
rect 165 -7 166 17
rect 170 -7 171 17
rect 165 -9 171 -7
rect 184 17 187 18
rect 184 13 185 17
rect 184 -9 187 13
<< ndcontact >>
rect 55 -26 59 -22
rect -23 -48 -19 -44
rect -4 -46 0 -42
rect 15 -48 19 -44
rect 48 -47 52 -43
rect 74 -46 78 -42
rect 112 -46 116 -42
rect 131 -26 135 -22
rect 138 -47 142 -43
rect 171 -48 175 -44
rect 190 -46 194 -42
rect 209 -48 213 -44
rect 55 -58 59 -54
rect 74 -57 78 -53
rect 93 -56 97 -52
rect 112 -57 116 -53
rect 131 -58 135 -54
<< pdcontact >>
rect 20 47 24 55
rect 39 30 43 34
rect 58 47 62 55
rect 128 47 132 55
rect 147 30 151 34
rect 166 47 170 54
rect 1 13 5 17
rect 20 -7 24 17
rect 39 13 43 17
rect 48 13 52 17
rect 55 3 59 7
rect 74 5 78 9
rect 93 -7 97 -3
rect 138 13 142 17
rect 112 5 116 9
rect 131 3 135 7
rect 147 13 151 17
rect 166 -7 170 17
rect 185 13 189 17
<< polysilicon >>
rect 25 57 26 58
rect 37 57 38 58
rect 25 56 38 57
rect 44 56 57 58
rect 133 56 146 58
rect 152 57 153 58
rect 164 57 165 58
rect 152 56 165 57
rect 25 27 38 29
rect 44 27 57 29
rect 133 27 146 29
rect 152 27 165 29
rect 6 19 7 20
rect 11 19 19 20
rect 6 18 19 19
rect 25 19 26 20
rect 48 22 51 23
rect 30 19 38 20
rect 25 18 38 19
rect 44 19 51 22
rect 79 19 83 20
rect 87 19 92 20
rect 44 18 47 19
rect 79 18 92 19
rect 98 19 103 20
rect 139 22 142 23
rect 107 19 111 20
rect 139 19 146 22
rect 98 18 111 19
rect 143 18 146 19
rect 152 19 160 20
rect 164 19 165 20
rect 152 18 165 19
rect 171 19 179 20
rect 183 19 184 20
rect 171 18 184 19
rect 60 10 61 11
rect 65 10 73 11
rect 60 9 73 10
rect 60 1 73 3
rect 117 10 125 11
rect 129 10 130 11
rect 117 9 130 10
rect 117 1 130 3
rect 6 -11 19 -9
rect 25 -11 38 -9
rect 44 -11 47 -9
rect 79 -11 92 -9
rect 98 -11 111 -9
rect 143 -11 146 -9
rect 152 -11 165 -9
rect 171 -11 184 -9
rect 60 -20 61 -19
rect 65 -20 73 -19
rect 60 -21 73 -20
rect 117 -20 125 -19
rect 129 -20 130 -19
rect 117 -21 130 -20
rect -18 -42 -5 -40
rect 1 -42 14 -40
rect 20 -44 47 -42
rect 20 -49 47 -47
rect 60 -49 73 -48
rect -18 -50 -5 -49
rect -18 -51 -17 -50
rect -13 -51 -5 -50
rect 1 -51 14 -49
rect 20 -51 73 -49
rect 1 -53 25 -51
rect 60 -52 73 -51
rect 79 -51 87 -50
rect 91 -51 92 -50
rect 79 -52 92 -51
rect 98 -51 99 -50
rect 176 -42 189 -40
rect 195 -42 208 -40
rect 143 -44 170 -42
rect 117 -49 130 -48
rect 143 -49 170 -47
rect 103 -51 111 -50
rect 98 -52 111 -51
rect 117 -51 170 -49
rect 176 -51 189 -49
rect 195 -50 208 -49
rect 195 -51 203 -50
rect 117 -52 130 -51
rect 165 -53 189 -51
rect 207 -51 208 -50
rect 60 -61 73 -59
rect 79 -61 92 -59
rect 98 -61 111 -59
rect 117 -61 130 -59
<< polycontact >>
rect 26 57 37 61
rect 153 57 164 61
rect 48 23 52 27
rect 138 23 142 27
rect 7 19 11 23
rect 26 19 30 23
rect 83 19 87 23
rect 103 19 107 23
rect 160 19 164 23
rect 179 19 183 23
rect 61 10 65 14
rect 125 10 129 14
rect 61 -20 65 -16
rect 125 -20 129 -16
rect -17 -54 -13 -50
rect 87 -51 91 -47
rect 99 -51 103 -47
rect 203 -54 207 -50
<< metal1 >>
rect -23 61 213 64
rect -23 57 26 61
rect 37 57 73 61
rect 77 57 113 61
rect 117 57 153 61
rect 164 57 213 61
rect -23 55 213 57
rect -23 47 20 55
rect 24 47 58 55
rect 62 47 128 55
rect 132 54 213 55
rect 132 47 166 54
rect 170 47 213 54
rect -23 46 213 47
rect -23 23 -10 27
rect 1 19 7 46
rect 20 19 26 23
rect 1 17 5 19
rect 20 17 24 19
rect 39 17 43 30
rect 56 23 134 27
rect 48 17 52 23
rect 20 -12 24 -7
rect -4 -16 20 -12
rect -4 -42 0 -16
rect 48 -43 52 13
rect 61 14 65 23
rect 125 14 129 23
rect 138 17 142 23
rect 147 17 151 30
rect 164 19 170 23
rect 183 19 189 46
rect 166 17 170 19
rect 55 -16 59 3
rect 55 -20 61 -16
rect 65 -19 84 -16
rect 65 -20 80 -19
rect 55 -22 59 -20
rect -23 -50 -19 -48
rect -23 -54 -17 -50
rect 15 -54 19 -48
rect 74 -53 78 -46
rect 93 -47 97 -7
rect 131 -16 135 3
rect 110 -19 125 -16
rect 114 -20 125 -19
rect 129 -20 135 -16
rect 131 -22 135 -20
rect 91 -51 99 -47
rect -23 -58 55 -54
rect 93 -52 97 -51
rect 112 -53 116 -46
rect 138 -43 142 13
rect 185 17 189 19
rect 166 -12 170 -7
rect 170 -16 213 -12
rect 190 -42 194 -16
rect 171 -54 175 -48
rect 209 -50 213 -48
rect 207 -54 213 -50
rect -23 -60 59 -58
rect 135 -58 213 -54
rect 131 -60 213 -58
rect -23 -71 213 -60
<< m2contact >>
rect 73 57 77 61
rect 113 57 117 61
rect -10 23 -6 27
rect 52 23 56 27
rect 134 23 138 27
rect 20 -16 24 -12
rect 74 9 78 13
rect 112 9 116 13
rect 80 -23 84 -19
rect 110 -23 114 -19
rect 166 -16 170 -12
<< metal2 >>
rect -6 23 52 27
rect 73 23 77 57
rect 113 23 117 57
rect 138 23 142 27
rect 74 13 78 23
rect 112 13 116 23
rect 24 -16 166 -12
rect 84 -23 110 -19
<< labels >>
rlabel metal1 4 60 4 60 5 Vdd
rlabel metal1 1 -58 1 -58 1 Gnd
rlabel metal2 110 -15 110 -15 7 Cascode
rlabel metal2 -4 25 -4 25 3 Bias
<< end >>
