magic
tech scmos
timestamp 1355110656
<< nwell >>
rect 216 -208 316 -207
rect 148 -297 316 -208
<< pwell >>
rect 148 -344 317 -297
<< ntransistor >>
rect 169 -313 172 -303
rect 178 -313 181 -303
rect 195 -313 198 -303
rect 201 -313 204 -303
rect 174 -338 177 -328
rect 192 -338 195 -328
rect 201 -338 204 -328
<< ptransistor >>
rect 174 -255 177 -235
rect 191 -255 194 -235
rect 204 -255 207 -235
rect 174 -289 177 -269
rect 183 -289 186 -269
rect 192 -289 195 -269
rect 201 -289 204 -269
<< ndiffusion >>
rect 168 -309 169 -303
rect 164 -313 169 -309
rect 172 -313 173 -303
rect 177 -313 178 -303
rect 181 -309 182 -303
rect 181 -313 186 -309
rect 194 -309 195 -303
rect 190 -313 195 -309
rect 198 -313 201 -303
rect 204 -313 205 -303
rect 169 -329 174 -328
rect 173 -333 174 -329
rect 169 -338 174 -333
rect 177 -329 183 -328
rect 177 -337 178 -329
rect 182 -337 183 -329
rect 177 -338 183 -337
rect 187 -329 192 -328
rect 191 -333 192 -329
rect 187 -338 192 -333
rect 195 -338 201 -328
rect 204 -329 209 -328
rect 204 -337 205 -329
rect 204 -338 209 -337
<< pdiffusion >>
rect 171 -236 174 -235
rect 173 -242 174 -236
rect 169 -246 174 -242
rect 173 -253 174 -246
rect 169 -254 174 -253
rect 171 -255 174 -254
rect 177 -236 182 -235
rect 177 -253 178 -236
rect 177 -255 182 -253
rect 186 -238 191 -235
rect 190 -242 191 -238
rect 186 -246 191 -242
rect 190 -253 191 -246
rect 186 -255 191 -253
rect 194 -241 204 -235
rect 194 -245 199 -241
rect 203 -245 204 -241
rect 194 -249 204 -245
rect 194 -253 199 -249
rect 203 -253 204 -249
rect 194 -255 204 -253
rect 207 -236 210 -235
rect 207 -253 208 -236
rect 207 -255 212 -253
rect 171 -270 174 -269
rect 173 -277 174 -270
rect 169 -281 174 -277
rect 173 -288 174 -281
rect 171 -289 174 -288
rect 177 -270 183 -269
rect 177 -288 178 -270
rect 182 -288 183 -270
rect 177 -289 183 -288
rect 186 -270 192 -269
rect 186 -277 187 -270
rect 191 -277 192 -270
rect 186 -281 192 -277
rect 186 -286 187 -281
rect 191 -286 192 -281
rect 186 -289 192 -286
rect 195 -270 201 -269
rect 195 -287 196 -270
rect 200 -287 201 -270
rect 195 -289 201 -287
rect 204 -270 207 -269
rect 204 -288 205 -270
rect 204 -289 207 -288
<< ndcontact >>
rect 164 -309 168 -303
rect 173 -313 177 -303
rect 182 -309 186 -303
rect 190 -309 194 -303
rect 205 -313 209 -303
rect 169 -333 173 -329
rect 178 -337 182 -329
rect 187 -333 191 -329
rect 205 -337 209 -329
<< pdcontact >>
rect 169 -242 173 -236
rect 169 -253 173 -246
rect 178 -253 182 -236
rect 186 -242 190 -238
rect 186 -253 190 -246
rect 199 -245 203 -241
rect 199 -253 203 -249
rect 208 -253 212 -236
rect 169 -277 173 -270
rect 169 -288 173 -281
rect 178 -288 182 -270
rect 187 -277 191 -270
rect 187 -286 191 -281
rect 196 -287 200 -270
rect 205 -288 209 -270
<< psubstratepdiff >>
rect 235 -332 239 -328
<< nsubstratendiff >>
rect 307 -221 311 -217
<< psubstratepcontact >>
rect 239 -332 243 -328
<< nsubstratencontact >>
rect 303 -221 307 -217
<< polysilicon >>
rect 174 -235 177 -233
rect 191 -235 194 -233
rect 204 -235 207 -233
rect 174 -269 177 -255
rect 191 -256 194 -255
rect 204 -256 207 -255
rect 181 -259 194 -256
rect 206 -260 207 -256
rect 194 -267 195 -263
rect 183 -269 186 -267
rect 192 -269 195 -267
rect 201 -269 204 -267
rect 174 -291 177 -289
rect 169 -294 177 -291
rect 169 -303 172 -294
rect 183 -297 186 -289
rect 178 -300 186 -297
rect 192 -298 195 -289
rect 178 -303 181 -300
rect 192 -301 198 -298
rect 195 -303 198 -301
rect 201 -303 204 -289
rect 169 -324 172 -313
rect 178 -316 181 -313
rect 195 -316 198 -313
rect 201 -315 204 -313
rect 180 -320 181 -316
rect 197 -320 198 -316
rect 185 -324 189 -322
rect 169 -327 177 -324
rect 185 -327 195 -324
rect 202 -326 203 -322
rect 174 -328 177 -327
rect 192 -328 195 -327
rect 201 -327 207 -326
rect 201 -328 204 -327
rect 174 -340 177 -338
rect 192 -340 195 -338
rect 201 -340 204 -338
<< polycontact >>
rect 181 -263 185 -259
rect 202 -260 206 -256
rect 190 -267 194 -263
rect 204 -299 208 -295
rect 176 -320 180 -316
rect 185 -322 189 -318
rect 193 -320 197 -316
rect 203 -326 207 -322
<< metal1 >>
rect 133 -199 334 -187
rect 134 -290 140 -199
rect 219 -211 305 -210
rect 218 -217 316 -211
rect 218 -221 303 -217
rect 307 -221 316 -217
rect 218 -232 316 -221
rect 179 -235 196 -232
rect 179 -236 182 -235
rect 193 -256 196 -235
rect 217 -244 221 -232
rect 212 -253 221 -244
rect 328 -251 334 -199
rect 191 -259 196 -256
rect 178 -263 181 -259
rect 191 -263 194 -259
rect 178 -270 182 -263
rect 199 -263 206 -260
rect 199 -270 202 -263
rect 200 -274 202 -270
rect 179 -289 182 -288
rect 134 -316 139 -290
rect 179 -292 186 -289
rect 182 -303 186 -292
rect 197 -303 200 -287
rect 209 -279 214 -253
rect 216 -303 219 -301
rect 134 -320 176 -316
rect 183 -318 186 -309
rect 197 -307 205 -303
rect 203 -313 205 -307
rect 212 -306 219 -303
rect 183 -322 185 -318
rect 197 -320 198 -316
rect 195 -337 198 -320
rect 203 -322 207 -313
rect 212 -316 216 -306
rect 210 -319 216 -316
rect 236 -317 311 -316
rect 210 -329 213 -319
rect 236 -324 316 -317
rect 209 -337 213 -329
rect 217 -328 316 -324
rect 217 -329 239 -328
rect 178 -340 198 -337
rect 221 -332 239 -329
rect 243 -332 316 -328
rect 221 -344 316 -332
<< m2contact >>
rect 213 -232 218 -211
rect 169 -246 173 -242
rect 186 -246 190 -242
rect 199 -241 203 -237
rect 199 -249 203 -245
rect 169 -281 173 -277
rect 187 -281 191 -277
rect 208 -299 212 -295
rect 216 -301 221 -297
rect 164 -313 168 -309
rect 190 -313 194 -309
rect 187 -329 191 -325
rect 169 -337 173 -333
rect 217 -344 221 -329
<< metal2 >>
rect 164 -232 213 -211
rect 164 -234 191 -232
rect 169 -242 191 -234
rect 173 -246 186 -242
rect 190 -246 191 -242
rect 169 -277 191 -246
rect 199 -244 203 -241
rect 199 -245 221 -244
rect 203 -249 221 -245
rect 173 -281 187 -277
rect 190 -299 208 -295
rect 216 -297 221 -249
rect 190 -301 194 -299
rect 143 -305 194 -301
rect 143 -349 151 -305
rect 168 -313 190 -309
rect 164 -325 194 -313
rect 164 -329 187 -325
rect 191 -329 194 -325
rect 164 -333 217 -329
rect 164 -337 169 -333
rect 173 -337 217 -333
rect 164 -344 217 -337
rect 332 -349 340 -313
rect 143 -356 340 -349
rect 143 -357 151 -356
<< labels >>
rlabel metal1 314 -344 316 -317 1 Vneg
rlabel nwell 315 -234 316 -211 1 Vpos
rlabel pwell 212 -344 214 -317 3 Vneg
rlabel metal2 219 -287 219 -287 1 D
rlabel metal1 138 -211 138 -211 3 Q
rlabel metal2 145 -331 145 -331 1 Qbar
rlabel polysilicon 170 -293 170 -293 1 T
rlabel metal1 180 -291 180 -291 1 N1
rlabel metal1 199 -293 199 -293 1 N2
<< end >>
