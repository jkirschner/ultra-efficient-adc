magic
tech scmos
timestamp 1355475848
<< nwell >>
rect -14 7 34 42
<< pwell >>
rect -14 -22 34 7
<< ntransistor >>
rect 2 -10 5 0
rect 11 -10 14 0
<< ptransistor >>
rect 2 15 5 35
rect 11 15 14 35
<< ndiffusion >>
rect -1 -7 2 0
rect 1 -10 2 -7
rect 5 -4 6 0
rect 10 -4 11 0
rect 5 -10 11 -4
rect 14 -7 17 0
rect 14 -10 15 -7
<< pdiffusion >>
rect -1 34 2 35
rect 1 30 2 34
rect -1 15 2 30
rect 5 15 11 35
rect 14 21 17 35
rect 14 17 15 21
rect 14 15 17 17
<< ndcontact >>
rect -3 -11 1 -7
rect 6 -4 10 0
rect 15 -11 19 -7
<< pdcontact >>
rect -3 30 1 34
rect 15 17 19 21
<< psubstratepcontact >>
rect 23 -15 27 -11
<< nsubstratencontact >>
rect 21 33 25 37
<< polysilicon >>
rect 2 35 5 37
rect 11 35 14 37
rect 2 7 5 15
rect 11 14 14 15
rect 2 0 5 3
rect 11 0 14 10
rect 2 -12 5 -10
rect 11 -12 14 -10
<< polycontact >>
rect 10 10 14 14
rect 1 3 5 7
<< metal1 >>
rect -14 37 34 42
rect -14 34 21 37
rect -14 30 -3 34
rect 1 33 21 34
rect 25 33 34 37
rect 1 30 34 33
rect -14 28 34 30
rect 19 17 21 21
rect -14 10 10 14
rect 17 11 21 17
rect 17 7 34 11
rect -14 3 1 7
rect 17 1 21 7
rect 8 0 21 1
rect 10 -4 21 0
rect -14 -11 -3 -7
rect 1 -11 15 -7
rect 19 -11 34 -7
rect -14 -15 23 -11
rect 27 -15 34 -11
rect -14 -22 34 -15
<< labels >>
rlabel metal1 -5 12 -5 12 3 A
rlabel metal1 -5 5 -5 5 3 B
rlabel metal1 19 8 19 8 7 Out
rlabel metal1 -10 32 -9 33 3 pos
rlabel metal1 -11 -11 -10 -10 3 neg
<< end >>
