magic
tech scmos
timestamp 1355237128
<< nwell >>
rect -27 53 141 95
rect 13 52 141 53
rect 13 51 124 52
rect 29 50 124 51
rect 39 49 112 50
<< pwell >>
rect -27 51 13 53
rect -27 50 29 51
rect 124 50 141 52
rect -27 49 39 50
rect 112 49 141 50
rect -27 8 141 49
rect 89 5 114 8
<< ntransistor >>
rect -15 29 -7 44
rect 0 44 2 47
rect 16 41 18 44
rect 24 34 26 37
rect 1 28 3 31
rect 36 28 44 43
rect 50 38 52 41
rect 66 38 69 41
rect 75 38 78 41
rect 92 38 94 41
rect 92 28 94 31
rect 102 28 104 31
rect 97 16 101 18
<< ptransistor >>
rect 4 73 6 79
rect 19 75 25 77
rect 0 60 2 66
rect 32 70 56 82
rect 67 76 83 82
rect 92 68 94 74
rect 100 68 102 74
rect 24 57 26 63
rect 32 57 35 61
rect 49 55 51 61
rect 66 55 69 61
rect 75 55 78 61
rect 92 55 94 61
<< ndiffusion >>
rect -16 29 -15 44
rect -7 41 -6 44
rect -2 44 0 47
rect 2 44 3 47
rect -2 41 -1 44
rect -7 39 -1 41
rect 15 41 16 44
rect 18 41 19 44
rect -7 31 -3 39
rect 31 37 36 43
rect 23 34 24 37
rect 26 34 27 37
rect -7 29 -6 31
rect 0 28 1 31
rect 3 28 4 31
rect 35 28 36 37
rect 44 41 49 43
rect 44 30 45 41
rect 49 38 50 41
rect 52 38 53 41
rect 65 38 66 41
rect 69 38 70 41
rect 74 38 75 41
rect 78 38 79 41
rect 91 38 92 41
rect 94 38 95 41
rect 44 28 49 30
rect 91 28 92 31
rect 94 28 95 31
rect 99 28 102 31
rect 104 30 110 31
rect 104 28 106 30
rect 97 18 101 19
rect 97 15 101 16
<< pdiffusion >>
rect 32 83 33 85
rect 43 83 47 87
rect 55 83 56 85
rect 32 82 56 83
rect 81 83 83 87
rect 67 82 83 83
rect 1 77 4 79
rect 3 73 4 77
rect 6 77 9 79
rect 19 78 21 80
rect 19 77 25 78
rect 6 73 7 77
rect -3 64 0 66
rect -1 60 0 64
rect 2 64 5 66
rect 2 60 3 64
rect 19 74 25 75
rect 23 72 25 74
rect 67 75 83 76
rect 32 69 56 70
rect 32 67 36 69
rect 49 67 56 69
rect 91 68 92 74
rect 94 70 95 74
rect 99 70 100 74
rect 94 68 100 70
rect 102 70 103 74
rect 102 68 105 70
rect 21 61 24 63
rect 23 57 24 61
rect 26 61 29 63
rect 26 57 27 61
rect 31 57 32 61
rect 35 57 36 61
rect 48 57 49 61
rect 46 55 49 57
rect 51 57 52 61
rect 51 55 54 57
rect 65 55 66 61
rect 69 59 75 61
rect 69 55 70 59
rect 74 55 75 59
rect 78 55 79 61
rect 91 55 92 61
rect 94 55 95 61
<< ndcontact >>
rect -20 29 -16 44
rect -6 41 -2 47
rect 3 43 7 47
rect 11 40 15 44
rect 19 41 23 45
rect 19 33 23 37
rect -6 27 0 31
rect 4 27 8 31
rect 27 28 35 37
rect 45 30 49 41
rect 53 37 57 41
rect 61 35 65 41
rect 70 37 74 41
rect 79 35 83 41
rect 87 36 91 41
rect 95 37 99 41
rect 87 26 91 31
rect 95 27 99 31
rect 106 26 110 30
rect 97 19 101 23
rect 97 11 101 15
<< pdcontact >>
rect 33 83 43 87
rect 47 83 55 87
rect 67 83 81 87
rect -1 73 3 77
rect 21 78 25 82
rect 7 73 11 77
rect -5 60 -1 64
rect 3 60 7 64
rect 19 70 23 74
rect 67 71 83 75
rect 36 65 49 69
rect 87 68 91 74
rect 95 70 99 74
rect 103 70 107 74
rect 19 57 23 61
rect 27 57 31 61
rect 36 57 40 61
rect 44 57 48 61
rect 52 57 56 61
rect 61 55 65 61
rect 70 55 74 59
rect 79 55 83 61
rect 87 55 91 61
rect 95 55 99 61
<< psubstratepdiff >>
rect 68 27 72 31
<< nsubstratendiff >>
rect -5 73 -1 77
<< psubstratepcontact >>
rect 64 27 68 31
<< nsubstratencontact >>
rect -9 73 -5 77
<< polysilicon >>
rect 4 79 6 81
rect 15 77 18 81
rect 15 75 19 77
rect 25 75 27 77
rect 4 71 6 73
rect 0 66 2 68
rect 0 47 2 60
rect -15 44 -7 46
rect 0 42 2 44
rect 15 46 18 75
rect 30 70 32 82
rect 56 73 58 82
rect 65 76 67 82
rect 83 78 84 82
rect 96 81 133 85
rect 83 76 85 78
rect 56 70 57 73
rect 92 74 94 81
rect 100 74 102 76
rect 92 66 94 68
rect 100 67 102 68
rect 24 63 26 65
rect 32 61 35 63
rect 49 61 51 63
rect 66 61 69 63
rect 75 61 78 63
rect 92 61 94 63
rect 16 44 18 46
rect 24 56 26 57
rect 16 39 18 41
rect 24 38 27 56
rect 32 55 35 57
rect 32 54 38 55
rect 32 52 34 54
rect 49 53 51 55
rect 49 48 52 53
rect 66 51 69 55
rect 75 51 78 55
rect 66 50 78 51
rect 92 50 94 55
rect 36 43 44 45
rect 67 46 77 50
rect 24 37 26 38
rect 1 31 3 34
rect -15 27 -7 29
rect 1 26 3 28
rect 24 29 26 34
rect 22 25 26 29
rect 50 41 52 44
rect 66 45 78 46
rect 66 41 69 45
rect 75 41 78 45
rect 92 41 94 46
rect 102 43 105 47
rect 50 36 52 38
rect 66 36 69 38
rect 75 36 78 38
rect 92 36 94 38
rect 92 31 94 33
rect 101 32 105 43
rect 102 31 104 32
rect 36 26 44 28
rect 92 23 94 28
rect 102 26 104 28
rect 126 18 133 81
rect 95 16 97 18
rect 101 16 133 18
<< polycontact >>
rect 3 81 7 85
rect 14 81 18 85
rect -4 51 0 55
rect 84 78 88 82
rect 92 81 96 85
rect 57 69 61 73
rect 99 63 103 67
rect 34 50 38 54
rect 48 44 52 48
rect 63 46 67 50
rect 77 46 81 50
rect 90 46 94 50
rect 1 34 5 38
rect -13 23 -9 27
rect 98 43 102 47
rect 22 21 26 25
rect 38 22 42 26
<< metal1 >>
rect 14 93 105 94
rect 14 91 110 93
rect 14 90 81 91
rect 91 90 110 91
rect 14 85 18 90
rect 55 83 67 87
rect 84 82 88 88
rect 25 78 29 82
rect 23 77 29 78
rect -5 68 -1 77
rect 11 73 14 74
rect 7 71 14 73
rect -20 51 -4 55
rect -20 44 -16 51
rect 3 47 7 60
rect 10 61 14 71
rect 26 70 29 77
rect 19 67 23 70
rect 19 64 31 67
rect 27 61 31 64
rect 10 57 19 61
rect 73 65 77 71
rect 103 74 110 90
rect 107 70 110 74
rect 36 61 40 65
rect 61 62 82 65
rect 61 61 65 62
rect 10 56 15 57
rect -6 35 -3 41
rect 1 40 7 43
rect 11 44 15 56
rect 27 48 31 57
rect 45 54 48 57
rect 79 61 82 62
rect 88 61 91 68
rect 95 61 103 63
rect 99 59 103 61
rect 99 55 101 59
rect 38 51 58 54
rect 55 50 58 51
rect 70 51 74 55
rect 1 38 5 40
rect 11 31 15 40
rect 19 47 31 48
rect 19 45 48 47
rect 23 44 48 45
rect 55 46 63 50
rect 97 50 101 55
rect 55 41 58 46
rect 70 41 74 47
rect 81 46 90 50
rect 97 47 117 50
rect 97 43 98 47
rect 102 43 117 47
rect 95 42 117 43
rect 95 41 101 42
rect 19 37 23 41
rect 8 27 15 31
rect 57 37 58 41
rect 61 34 65 35
rect 79 34 83 35
rect 49 30 51 34
rect 45 27 51 30
rect 55 31 79 34
rect 55 27 64 31
rect 68 27 79 31
rect 99 37 101 41
rect 87 31 91 36
rect -9 23 22 24
rect -13 21 22 23
rect 22 16 26 21
rect 38 20 42 22
rect 97 23 101 27
rect 113 16 117 42
rect 22 15 94 16
rect 103 15 117 16
rect 22 12 97 15
rect 94 11 97 12
rect 101 13 117 15
rect 101 12 115 13
rect 101 11 103 12
<< m2contact >>
rect 7 81 11 85
rect 43 83 47 87
rect -5 64 -1 68
rect 3 64 7 68
rect 29 70 33 74
rect 57 73 61 77
rect 95 74 99 78
rect 52 61 56 65
rect 106 66 110 70
rect -6 31 -2 35
rect 70 47 74 51
rect 31 37 35 41
rect 51 27 55 34
rect 79 27 83 34
rect 99 27 103 31
rect 106 30 110 34
<< metal2 >>
rect 3 68 7 85
rect 14 83 43 87
rect 47 83 99 87
rect 14 80 99 83
rect 14 79 53 80
rect 14 78 20 79
rect -5 60 -1 64
rect 10 60 20 78
rect 29 66 35 70
rect -5 55 20 60
rect 31 41 35 66
rect 43 67 53 79
rect 95 78 99 80
rect 61 73 65 74
rect 57 70 65 73
rect 43 65 56 67
rect 43 61 52 65
rect 43 57 56 61
rect 61 59 65 70
rect 106 61 110 66
rect 61 55 74 59
rect 70 51 74 55
rect 106 53 115 61
rect 106 34 110 53
rect -2 31 51 34
rect -6 27 51 31
rect 83 31 103 34
rect 83 27 99 31
<< labels >>
rlabel metal1 -11 22 -11 22 1 Out
rlabel metal1 40 21 40 21 1 Vpw1
rlabel metal1 86 87 86 87 6 Vpw2
rlabel metal2 108 50 108 50 7 OutB
rlabel metal1 99 50 99 50 1 Out
rlabel polysilicon 129 22 129 22 7 Reset
rlabel polysilicon 93 24 93 24 1 ResetB
rlabel polysilicon 25 30 25 30 1 Out
rlabel ndcontact 47 30 47 30 7 Vneg
<< end >>
