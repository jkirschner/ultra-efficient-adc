magic
tech scmos
timestamp 1355674183
<< metal1 >>
rect 353 3040 358 3047
rect 353 2900 358 2907
rect -787 2604 -48 2619
rect 169 2592 222 2597
rect 356 2582 360 2584
rect 334 2514 360 2582
rect 377 2522 381 2582
rect 386 2531 391 2581
rect 386 2525 463 2531
rect 377 2517 436 2522
rect 334 2511 410 2514
rect -874 2188 -843 2230
rect -8 1597 10 2507
rect 335 2494 410 2511
rect 177 1953 185 2133
rect 418 1563 436 2517
rect 406 1554 436 1563
rect 445 1606 463 2525
rect 406 1529 414 1554
rect 445 1532 462 1606
rect 361 1503 366 1512
rect 445 1511 463 1532
rect -2597 1005 -2585 1021
rect 19 -9 37 19
rect 48 0 79 7
rect 48 -8 52 0
rect 129 -7 152 16
rect 65 -17 152 -7
rect 47 -75 51 -52
<< m2contact >>
rect -798 2604 -787 2619
rect 222 2590 230 2597
rect 18 2580 45 2587
rect 19 2504 46 2511
rect 177 2133 185 2140
rect 445 1499 463 1511
<< metal2 >>
rect -392 2510 -386 2625
rect -107 2569 -101 2625
rect -107 2564 -62 2569
rect 18 2511 45 2580
rect -392 2497 -62 2510
rect 18 2504 19 2511
rect 158 2509 164 2581
rect 179 2514 184 2582
rect 171 2509 184 2514
rect 222 2140 230 2590
rect 185 2133 230 2140
rect 378 1511 463 1512
rect 378 1499 445 1511
use stateMachine  stateMachine_0
timestamp 1355540337
transform 1 0 -1265 0 1 3050
box -14 -441 1196 68
use msb_registers  msb_registers_0
timestamp 1355455137
transform 0 1 227 1 0 2875
box -295 -224 301 222
use Comparator  Comparator_0
timestamp 1355605154
transform 0 1 -1060 1 0 1639
box -6 -28 815 195
use lsb_registers_Layout  lsb_registers_Layout_0
timestamp 1355599904
transform 0 1 263 -1 0 1521
box -990 -263 1521 160
use NOT  NOT_0
timestamp 1355475633
transform 0 1 42 -1 0 -12
box -5 -23 43 41
<< labels >>
rlabel metal1 49 -72 49 -72 1 GO?
<< end >>
