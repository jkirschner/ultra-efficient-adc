* SPICE3 file created from Comparator.ext - technology: scmos

.subckt GainLatch_layout PosA PosD Disable Vm Vp Dout Vneg Vbias Cascode
M1000 a_26_61# Cascode N1 PosA pfet w=4.8u l=2.4u
+ ad=29.52p pd=43.2u as=27p ps=46.8u 
M1001 PosA Vbias a_26_61# PosA pfet w=9u l=18u
+ ad=16.2p pd=21.6u as=0p ps=0u 
M1002 a_26_61# Vbias PosA PosA pfet w=9u l=18u
+ ad=0p pd=0u as=0p ps=0u 
M1003 N1 Cascode a_26_61# PosA pfet w=4.8u l=2.4u
+ ad=0p pd=0u as=0p ps=0u 
M1004 PosD Disable a_19_27# PosA pfet w=4.5u l=2.7u
+ ad=16.2p pd=25.2u as=15.48p ps=34.8u 
M1005 a_33_11# a_33_11# PosD PosA pfet w=4.5u l=2.7u
+ ad=13.5p pd=24u as=0p ps=0u 
M1006 N1 Vp N3 PosA pfet w=3.6u l=3.6u
+ ad=0p pd=0u as=10.8p ps=20.4u 
M1007 N2 a_80_23# N1 PosA pfet w=3.6u l=3.6u
+ ad=6.48p pd=10.8u as=0p ps=0u 
M1008 N1 a_80_23# N2 PosA pfet w=3.6u l=3.6u
+ ad=0p pd=0u as=0p ps=0u 
M1009 N3 Vp N1 PosA pfet w=3.6u l=3.6u
+ ad=0p pd=0u as=0p ps=0u 
M1010 PosD a_33_11# a_33_11# PosA pfet w=4.5u l=2.7u
+ ad=0p pd=0u as=0p ps=0u 
M1011 a_19_27# Disable PosD PosA pfet w=4.5u l=2.7u
+ ad=0p pd=0u as=0p ps=0u 
M1012 Dout a_33_11# a_19_27# PosA pfet w=0.9u l=0.6u
+ ad=3.42p pd=10.8u as=0p ps=0u 
M1013 a_19_27# a_33_11# Dout PosA pfet w=0.9u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1014 Dout Disable Vneg Vneg nfet w=3.6u l=1.8u
+ ad=16.92p pd=36u as=36.72p ps=74.4u 
M1015 Vneg N3 Dout Vneg nfet w=2.4u l=2.7u
+ ad=0p pd=0u as=0p ps=0u 
M1016 N3 N3 Vneg Vneg nfet w=2.4u l=2.7u
+ ad=4.32p pd=8.4u as=0p ps=0u 
M1017 Vneg N3 N3 Vneg nfet w=2.4u l=2.7u
+ ad=0p pd=0u as=0p ps=0u 
M1018 Dout N3 Vneg Vneg nfet w=2.4u l=2.7u
+ ad=0p pd=0u as=0p ps=0u 
M1019 Vneg Disable Dout Vneg nfet w=3.6u l=1.8u
+ ad=0p pd=0u as=0p ps=0u 
M1020 a_33_11# Dout Vneg Vneg nfet w=3.6u l=1.8u
+ ad=16.92p pd=36u as=0p ps=0u 
M1021 Vneg N2 a_33_11# Vneg nfet w=2.4u l=2.7u
+ ad=0p pd=0u as=0p ps=0u 
M1022 N2 N2 Vneg Vneg nfet w=2.4u l=2.7u
+ ad=4.32p pd=8.4u as=0p ps=0u 
M1023 Vneg N2 N2 Vneg nfet w=2.4u l=2.7u
+ ad=0p pd=0u as=0p ps=0u 
M1024 a_33_11# N2 Vneg Vneg nfet w=2.4u l=2.7u
+ ad=0p pd=0u as=0p ps=0u 
M1025 Vneg Dout a_33_11# Vneg nfet w=3.6u l=1.8u
+ ad=0p pd=0u as=0p ps=0u 
.ends

.subckt doublePreamp PosA V+ Thresh V- Bias Vneg Input Cascode
** SOURCE/DRAIN TIED
M1000 PosA PosA PosA PosA pfet w=1.8u l=0.9u
+ ad=34.2p pd=73.2u as=0p ps=0u 
M1001 a_32_49# Bias PosA PosA pfet w=8.1u l=3.9u
+ ad=17.82p pd=39.6u as=0p ps=0u 
M1002 a_24_22# Cascode a_32_49# PosA pfet w=1.8u l=0.9u
+ ad=12.78p pd=30u as=0p ps=0u 
M1003 a_32_49# Cascode a_24_22# PosA pfet w=1.8u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1004 PosA Bias a_32_49# PosA pfet w=8.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
** SOURCE/DRAIN TIED
M1005 PosA PosA PosA PosA pfet w=1.8u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1006 V- PosA PosA PosA pfet w=1.5u l=0.9u
+ ad=13.5p pd=24u as=0p ps=0u 
M1007 a_24_22# Input V- PosA pfet w=1.5u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1008 V+ Thresh a_24_22# PosA pfet w=1.5u l=0.9u
+ ad=4.14p pd=12u as=0p ps=0u 
M1009 a_24_22# Thresh V+ PosA pfet w=1.5u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1010 V- Input a_24_22# PosA pfet w=1.5u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1011 PosA PosA V- PosA pfet w=1.5u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1012 V- Vneg Vneg Vneg nfet w=1.5u l=0.9u
+ ad=5.4p pd=13.2u as=12.24p ps=28.8u 
M1013 Vneg V- V- Vneg nfet w=1.5u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1014 V+ V- Vneg Vneg nfet w=1.5u l=0.9u
+ ad=4.14p pd=12u as=0p ps=0u 
M1015 Vneg V- V+ Vneg nfet w=1.5u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1016 V- V- Vneg Vneg nfet w=1.5u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1017 Vneg Vneg V- Vneg nfet w=1.5u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
.ends

.subckt doubleBiasGen PosA Bias Vneg Cascode
M1000 a_38_n9# PosA PosA PosA pfet w=8.1u l=3.9u
+ ad=29.16p pd=39.6u as=68.58p ps=154.8u 
M1001 PosA Bias a_38_n9# PosA pfet w=8.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1002 a_146_n9# Bias PosA PosA pfet w=8.1u l=3.9u
+ ad=29.16p pd=39.6u as=0p ps=0u 
M1003 PosA PosA a_146_n9# PosA pfet w=8.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1004 Cascode PosA PosA PosA pfet w=8.1u l=3.9u
+ ad=29.16p pd=39.6u as=0p ps=0u 
M1005 a_38_n9# Cascode Cascode PosA pfet w=8.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1006 Bias Bias a_38_n9# PosA pfet w=8.1u l=0.9u
+ ad=16.02p pd=38.4u as=0p ps=0u 
M1007 PosA Bias a_1_n53# PosA pfet w=1.8u l=3.9u
+ ad=0p pd=0u as=4.68p ps=13.2u 
M1008 a_79_n61# Bias PosA PosA pfet w=8.1u l=3.9u
+ ad=14.58p pd=19.8u as=0p ps=0u 
M1009 PosA Bias a_79_n61# PosA pfet w=8.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1010 a_1_n53# Bias PosA PosA pfet w=1.8u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1011 a_146_n9# Bias Bias PosA pfet w=8.1u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1012 Cascode Cascode a_146_n9# PosA pfet w=8.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1013 PosA PosA Cascode PosA pfet w=8.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1014 Cascode Vneg Vneg Vneg nfet w=2.1u l=3.9u
+ ad=7.56p pd=15.6u as=16.2p ps=44.4u 
M1015 Vneg a_1_n53# Cascode Vneg nfet w=2.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1016 Bias a_1_n53# Vneg Vneg nfet w=0.9u l=8.1u
+ ad=3.42p pd=10.8u as=0p ps=0u 
M1017 a_73_n59# a_1_n53# a_1_n53# Vneg nfet w=8.1u l=3.9u
+ ad=11.79p pd=27u as=16.02p ps=38.4u 
M1018 a_1_n53# a_1_n53# a_111_n59# Vneg nfet w=8.1u l=3.9u
+ ad=0p pd=0u as=11.79p ps=27u 
M1019 Vneg a_1_n53# Bias Vneg nfet w=0.9u l=8.1u
+ ad=0p pd=0u as=0p ps=0u 
M1020 Cascode a_1_n53# Vneg Vneg nfet w=2.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1021 Vneg Vneg Cascode Vneg nfet w=2.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1022 a_73_n59# a_1_n53# Vneg Vneg nfet w=2.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1023 a_79_n61# a_79_n61# a_73_n59# Vneg nfet w=2.1u l=3.9u
+ ad=3.78p pd=7.8u as=0p ps=0u 
M1024 a_111_n59# a_79_n61# a_79_n61# Vneg nfet w=2.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1025 Vneg a_1_n53# a_111_n59# Vneg nfet w=2.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
.ends


* Top level circuit Comparator

XGainLatch_layout_0 doublePreamp_0/PosA PosD Disable doublePreamp_0/V- doublePreamp_0/V+ Out doublePreamp_0/Vneg Bias doublePreamp_0/Cascode GainLatch_layout
XdoublePreamp_0 doublePreamp_0/PosA doublePreamp_0/V+ Thresh doublePreamp_0/V- Bias doublePreamp_0/Vneg Input doublePreamp_0/Cascode doublePreamp
XdoubleBiasGen_0 doublePreamp_0/PosA Bias doublePreamp_0/Vneg doublePreamp_0/Cascode doubleBiasGen
.end

