magic
tech scmos
timestamp 1355476235
<< nwell >>
rect 38 27 105 68
<< pwell >>
rect 38 1 105 27
<< ntransistor >>
rect 62 11 65 21
rect 79 11 82 21
rect 88 11 91 21
<< ptransistor >>
rect 62 33 65 53
rect 79 33 82 53
rect 88 33 91 53
<< ndiffusion >>
rect 59 16 62 21
rect 61 12 62 16
rect 59 11 62 12
rect 65 20 68 21
rect 65 16 66 20
rect 76 16 79 21
rect 65 11 68 16
rect 78 12 79 16
rect 76 11 79 12
rect 82 16 88 21
rect 82 12 83 16
rect 87 12 88 16
rect 82 11 88 12
rect 91 20 94 21
rect 91 16 92 20
rect 91 11 94 16
<< pdiffusion >>
rect 59 52 62 53
rect 61 48 62 52
rect 59 33 62 48
rect 65 38 68 53
rect 76 46 79 53
rect 78 42 79 46
rect 65 34 66 38
rect 65 33 68 34
rect 76 33 79 42
rect 82 39 88 53
rect 82 35 83 39
rect 87 35 88 39
rect 82 33 88 35
rect 91 49 92 53
rect 91 33 94 49
<< ndcontact >>
rect 57 12 61 16
rect 66 16 70 20
rect 74 12 78 16
rect 83 12 87 16
rect 92 16 96 20
<< pdcontact >>
rect 57 48 61 52
rect 74 42 78 46
rect 66 34 70 38
rect 83 35 87 39
rect 92 49 96 53
<< psubstratepcontact >>
rect 98 4 102 8
<< nsubstratencontact >>
rect 69 61 73 65
<< polysilicon >>
rect 62 54 82 56
rect 62 53 65 54
rect 79 53 82 54
rect 88 53 91 55
rect 62 29 65 33
rect 63 25 65 29
rect 62 21 65 25
rect 79 21 82 33
rect 88 28 91 33
rect 88 21 91 24
rect 62 9 65 11
rect 79 9 82 11
rect 88 9 91 11
<< polycontact >>
rect 59 25 63 29
rect 87 24 91 28
<< metal1 >>
rect 38 65 105 68
rect 38 61 69 65
rect 73 61 105 65
rect 38 57 105 61
rect 57 52 61 57
rect 74 49 92 53
rect 38 39 42 43
rect 78 42 98 46
rect 38 32 49 36
rect 38 25 59 29
rect 66 28 70 34
rect 66 24 87 28
rect 66 20 70 24
rect 94 21 98 42
rect 92 20 98 21
rect 96 16 98 20
rect 57 9 61 12
rect 38 8 105 9
rect 38 4 98 8
rect 102 4 105 8
rect 38 1 105 4
<< m2contact >>
rect 70 49 74 53
rect 42 39 46 43
rect 74 38 78 42
rect 49 32 53 36
rect 83 31 87 35
rect 101 29 105 33
rect 74 16 78 20
rect 83 16 87 20
<< metal2 >>
rect 64 49 70 53
rect 64 44 68 49
rect 42 43 68 44
rect 46 39 68 43
rect 42 24 46 39
rect 74 34 78 38
rect 53 32 78 34
rect 49 30 78 32
rect 87 31 101 33
rect 83 29 101 31
rect 42 20 78 24
rect 83 20 87 29
<< labels >>
rlabel m2contact 103 31 103 31 7 Out
rlabel metal1 59 58 59 58 5 Vdd
rlabel metal1 58 7 58 7 1 Gnd
rlabel metal1 50 27 50 27 1 S
rlabel metal1 39 41 39 41 3 In1
rlabel metal1 39 34 39 34 3 In2
<< end >>
