magic
tech scmos
timestamp 1355429379
<< ntransistor >>
rect 2 -10 5 0
rect 11 -10 14 0
<< ptransistor >>
rect 2 15 5 35
rect 11 15 14 35
<< ndiffusion >>
rect -1 -7 2 0
rect 1 -10 2 -7
rect 5 -4 6 0
rect 10 -4 11 0
rect 5 -10 11 -4
rect 14 -7 17 0
rect 14 -10 15 -7
<< pdiffusion >>
rect -1 34 2 35
rect 1 30 2 34
rect -1 15 2 30
rect 5 15 11 35
rect 14 21 17 35
rect 14 17 15 21
rect 14 15 17 17
<< ndcontact >>
rect -3 -11 1 -7
rect 6 -4 10 0
rect 15 -11 19 -7
<< pdcontact >>
rect -3 30 1 34
rect 15 17 19 21
<< polysilicon >>
rect 2 35 5 37
rect 11 35 14 37
rect 2 7 5 15
rect 11 14 14 15
rect 2 0 5 3
rect 11 0 14 10
rect 2 -12 5 -10
rect 11 -12 14 -10
<< polycontact >>
rect 10 10 14 14
rect 1 3 5 7
<< metal1 >>
rect -7 34 25 37
rect -7 30 -3 34
rect 1 30 25 34
rect -7 28 25 30
rect 19 17 21 21
rect -7 10 10 14
rect 17 10 21 17
rect 17 7 25 10
rect -7 3 1 7
rect 17 1 21 7
rect 8 0 21 1
rect 10 -4 21 0
rect -7 -11 -3 -7
rect 1 -11 15 -7
rect 19 -11 25 -7
rect -7 -15 25 -11
<< labels >>
rlabel metal1 7 -14 7 -14 1 Gnd
rlabel metal1 -5 35 -5 35 4 Vdd
rlabel metal1 -5 12 -5 12 3 A
rlabel metal1 -5 5 -5 5 3 B
rlabel metal1 19 8 19 8 7 Out
<< end >>
