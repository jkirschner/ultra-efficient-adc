magic
tech scmos
timestamp 1355639073
<< nwell >>
rect -531 1412 -521 1420
<< pwell >>
rect -529 1306 -525 1309
rect -529 1290 -525 1293
<< metal1 >>
rect -787 2604 -48 2619
rect -28 2604 -6 2619
rect -874 2188 -843 2230
rect -19 1600 8 2524
rect 19 2510 45 2532
rect 87 2524 174 2532
rect 192 2518 197 2525
rect 154 2513 197 2518
rect 335 2526 372 2532
rect 335 2511 360 2526
rect 386 2522 390 2533
rect 403 2527 461 2533
rect 386 2514 436 2522
rect 69 2496 75 2497
rect 335 2493 410 2511
rect 419 1554 436 2514
rect 378 1544 436 1554
rect 378 1534 386 1544
rect 444 1536 461 2527
rect 409 1527 461 1536
rect -531 1412 -521 1420
rect -529 1306 -525 1309
rect -529 1290 -525 1293
rect -2597 1005 -2585 1021
<< m2contact >>
rect -798 2604 -787 2619
rect -6 2604 8 2619
rect -19 2524 8 2532
rect 81 2524 87 2532
rect 192 2525 197 2533
rect 147 2513 154 2519
rect 377 2527 381 2533
rect 399 2527 403 2533
rect 69 2497 75 2510
<< metal2 >>
rect -392 2510 -386 2625
rect -107 2569 -101 2625
rect -6 2619 9 2620
rect 8 2604 9 2619
rect -107 2564 -62 2569
rect -20 2564 154 2569
rect 8 2524 81 2532
rect 147 2519 154 2564
rect 158 2510 164 2532
rect 179 2515 184 2532
rect 197 2527 377 2533
rect 381 2527 399 2533
rect 197 2525 403 2527
rect 171 2510 184 2515
rect -392 2497 -62 2510
rect -20 2497 69 2510
use stateMachine  stateMachine_0
timestamp 1355540337
transform 1 0 -1265 0 1 3050
box -14 -441 1196 68
use msb_registers  msb_registers_0
timestamp 1355455137
transform 0 1 227 1 0 2825
box -295 -224 301 222
use Comparator  Comparator_0
timestamp 1355605154
transform 0 1 -1060 1 0 1639
box -6 -28 815 195
use AnalogSwitch  AnalogSwitch_0
timestamp 1355620377
transform 1 0 -686 0 1 1376
box -325 -461 424 47
use lsb_registers_Layout  lsb_registers_Layout_0
timestamp 1355599904
transform 0 1 263 -1 0 1521
box -990 -263 1521 160
<< end >>
