* SPICE3 file created from AnalogSwitch.ext - technology: scmos

M1000 CLC1 NOT_0/In pos pos pfet w=6u l=0.9u
+ ad=6.12p pd=15u as=186.84p ps=264u 
M1001 CLC1 NOT_0/In neg neg nfet w=3u l=0.9u
+ ad=3.42p pd=9u as=79.74p ps=202.8u 
M1002 NOR_0/a_5_15# NOR_0/B pos pos pfet w=6u l=0.9u
+ ad=10.8p pd=15.6u as=0p ps=0u 
M1003 NOT_0/In RST_IR NOR_0/a_5_15# pos pfet w=6u l=0.9u
+ ad=6.12p pd=15u as=0p ps=0u 
M1004 NOT_0/In NOR_0/B neg neg nfet w=3u l=0.9u
+ ad=5.4p pd=9.6u as=0p ps=0u 
M1005 neg RST_IR NOT_0/In neg nfet w=3u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1006 NOR_2/a_5_15# NOR_2/B pos pos pfet w=6u l=0.9u
+ ad=10.8p pd=15.6u as=0p ps=0u 
M1007 NOR_0/B COb NOR_2/a_5_15# pos pfet w=6u l=0.9u
+ ad=6.12p pd=15u as=0p ps=0u 
M1008 NOR_0/B NOR_2/B neg neg nfet w=3u l=0.9u
+ ad=5.4p pd=9.6u as=0p ps=0u 
M1009 neg COb NOR_0/B neg nfet w=3u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1010 NOR_2/B RST_C1_CO? pos pos pfet w=6u l=0.9u
+ ad=6.12p pd=15u as=0p ps=0u 
M1011 NOR_2/B RST_C1_CO? neg neg nfet w=3u l=0.9u
+ ad=3.42p pd=9u as=0p ps=0u 
M1012 CLC2 NOT_1/In pos pos pfet w=6u l=0.9u
+ ad=6.12p pd=15u as=0p ps=0u 
M1013 CLC2 NOT_1/In neg neg nfet w=3u l=0.9u
+ ad=3.42p pd=9u as=0p ps=0u 
M1014 NOR_1/a_5_15# RST_IR pos pos pfet w=6u l=0.9u
+ ad=10.8p pd=15.6u as=0p ps=0u 
M1015 NOT_1/In NOR_1/A NOR_1/a_5_15# pos pfet w=6u l=0.9u
+ ad=6.12p pd=15u as=0p ps=0u 
M1016 NOT_1/In RST_IR neg neg nfet w=3u l=0.9u
+ ad=5.4p pd=9.6u as=0p ps=0u 
M1017 neg NOR_1/A NOT_1/In neg nfet w=3u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1018 NOR_3/a_5_15# COb pos pos pfet w=6u l=0.9u
+ ad=10.8p pd=15.6u as=0p ps=0u 
M1019 NOR_1/A NOR_3/A NOR_3/a_5_15# pos pfet w=6u l=0.9u
+ ad=6.12p pd=15u as=0p ps=0u 
M1020 NOR_1/A COb neg neg nfet w=3u l=0.9u
+ ad=5.4p pd=9.6u as=0p ps=0u 
M1021 neg NOR_3/A NOR_1/A neg nfet w=3u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1022 NOR_3/A RST_C2_CO? pos pos pfet w=6u l=0.9u
+ ad=6.12p pd=15u as=0p ps=0u 
M1023 NOR_3/A RST_C2_CO? neg neg nfet w=3u l=0.9u
+ ad=3.42p pd=9u as=0p ps=0u 
M1024 a_n13_n17# Iin? pos pos pfet w=6u l=0.9u
+ ad=10.8p pd=15.6u as=0p ps=0u 
M1025 pos C1? a_n13_n17# pos pfet w=6u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1026 a_n1_n33# C2? pos pos pfet w=6u l=0.9u
+ ad=10.8p pd=15.6u as=0p ps=0u 
M1027 pos Iin? a_n1_n33# pos pfet w=6u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1028 a_15_n33# a_n13_n17# pos pos pfet w=6u l=0.9u
+ ad=10.8p pd=15.6u as=0p ps=0u 
M1029 pos a_n1_n33# a_15_n33# pos pfet w=6u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1030 a_64_n23# Iin? pos pos pfet w=6u l=0.9u
+ ad=6.48p pd=15u as=0p ps=0u 
M1031 a_77_n33# a_64_n23# pos pos pfet w=6u l=0.9u
+ ad=10.8p pd=15.6u as=0p ps=0u 
M1032 pos C1? a_77_n33# pos pfet w=6u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1033 a_88_n33# a_64_n23# pos pos pfet w=6u l=0.9u
+ ad=10.8p pd=15.6u as=0p ps=0u 
M1034 pos C2? a_88_n33# pos pfet w=6u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1035 a_112_n33# a_88_n33# pos pos pfet w=6u l=0.9u
+ ad=10.8p pd=15.6u as=0p ps=0u 
M1036 pos a_77_n33# a_112_n33# pos pfet w=6u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1037 a_n5_n23# Iin? a_n13_n17# neg nfet w=3u l=0.9u
+ ad=5.4p pd=9.6u as=3.42p ps=9u 
M1038 neg C1? a_n5_n23# neg nfet w=3u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1039 a_13_n23# C2? neg neg nfet w=3u l=0.9u
+ ad=5.4p pd=9.6u as=0p ps=0u 
M1040 a_n1_n33# Iin? a_13_n23# neg nfet w=3u l=0.9u
+ ad=4.5p pd=9u as=0p ps=0u 
M1041 a_39_n23# a_n13_n17# neg neg nfet w=3u l=0.9u
+ ad=3.6p pd=8.4u as=0p ps=0u 
M1042 a_15_n33# a_n1_n33# a_39_n23# neg nfet w=3u l=0.9u
+ ad=4.41p pd=9u as=0p ps=0u 
M1043 a_64_n23# Iin? neg neg nfet w=3u l=0.9u
+ ad=3.42p pd=9u as=0p ps=0u 
M1044 a_81_n23# a_64_n23# neg neg nfet w=3u l=0.9u
+ ad=5.4p pd=9.6u as=0p ps=0u 
M1045 a_77_n33# C1? a_81_n23# neg nfet w=3u l=0.9u
+ ad=3.42p pd=9u as=0p ps=0u 
M1046 a_107_n23# a_64_n23# neg neg nfet w=3u l=0.9u
+ ad=5.4p pd=9.6u as=0p ps=0u 
M1047 a_88_n33# C2? a_107_n23# neg nfet w=3u l=0.9u
+ ad=3.42p pd=9u as=0p ps=0u 
M1048 a_133_n23# a_88_n33# neg neg nfet w=3u l=0.9u
+ ad=5.4p pd=9.6u as=0p ps=0u 
M1049 a_112_n33# a_77_n33# a_133_n23# neg nfet w=3u l=0.9u
+ ad=3.42p pd=9u as=0p ps=0u 
M1050 Iin a_n13_n17# VC1 pos pfet w=1.8u l=0.6u
+ ad=5.58p pd=13.8u as=4.68p ps=13.2u 
M1051 VC2 a_n1_n33# Iin pos pfet w=1.8u l=0.6u
+ ad=5.04p pd=13.2u as=0p ps=0u 
M1052 neg a_15_n33# Iin pos pfet w=1.8u l=0.6u
+ ad=17.64p pd=56.4u as=0p ps=0u 
M1053 Iref a_77_n33# VC1 pos pfet w=1.8u l=0.6u
+ ad=7.2p pd=15.6u as=0p ps=0u 
M1054 VC2 a_88_n33# Iref pos pfet w=1.8u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1055 neg a_112_n33# Iref pos pfet w=1.8u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1056 VC1 CLC1 neg neg nfet w=7.2u l=0.6u
+ ad=7.2p pd=17.4u as=0p ps=0u 
M1057 VC2 CLC2 neg neg nfet w=7.2u l=0.6u
+ ad=7.2p pd=17.4u as=0p ps=0u 
C0 neg VC1 10033.7fF
C1 neg VC2 10030.9fF
