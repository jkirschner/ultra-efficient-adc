magic
tech scmos
timestamp 1355075313
<< ntransistor >>
rect -38 27 -36 39
rect -38 2 -35 12
rect -8 -23 -5 -13
rect 1 -23 4 -13
rect 10 -23 13 -13
rect 19 -23 22 -13
rect 36 -23 39 -13
rect 43 -23 46 -13
rect 61 -23 64 -13
rect 78 -23 81 -13
rect 87 -23 90 -13
rect 104 -23 107 -13
rect 113 -23 116 -13
rect 130 -23 133 -13
rect 139 -23 142 -13
<< ptransistor >>
rect -59 31 -57 35
rect -59 1 -56 21
rect -8 -1 -5 19
rect 1 -1 4 19
rect 10 -1 13 19
rect 19 -1 22 19
rect 28 -1 31 19
rect 37 -1 40 19
rect 61 -1 64 19
rect 78 -1 81 19
rect 87 -1 90 19
rect 104 -1 107 19
rect 113 -1 116 19
rect 130 -1 133 19
rect 139 -1 142 19
<< ndiffusion >>
rect -41 27 -38 39
rect -36 27 -33 39
rect -41 2 -38 12
rect -35 2 -32 12
rect -9 -17 -8 -13
rect -11 -23 -8 -17
rect -5 -23 1 -13
rect 4 -20 10 -13
rect 4 -23 5 -20
rect 9 -23 10 -20
rect 13 -23 19 -13
rect 22 -17 23 -13
rect 22 -23 27 -17
rect 33 -19 36 -13
rect 35 -23 36 -19
rect 39 -23 43 -13
rect 46 -17 47 -13
rect 46 -23 51 -17
rect 58 -19 61 -13
rect 60 -23 61 -19
rect 64 -17 65 -13
rect 64 -23 67 -17
rect 75 -19 78 -13
rect 77 -23 78 -19
rect 81 -23 87 -13
rect 90 -17 91 -13
rect 90 -23 93 -17
rect 101 -19 104 -13
rect 103 -23 104 -19
rect 107 -23 113 -13
rect 116 -17 117 -13
rect 116 -23 119 -17
rect 127 -19 130 -13
rect 129 -23 130 -19
rect 133 -23 139 -13
rect 142 -17 143 -13
rect 142 -23 145 -17
<< pdiffusion >>
rect -62 31 -59 35
rect -57 31 -54 35
rect -62 1 -59 21
rect -56 1 -53 21
rect -11 17 -8 19
rect -9 13 -8 17
rect -11 -1 -8 13
rect -5 5 1 19
rect -5 1 -4 5
rect 0 1 1 5
rect -5 -1 1 1
rect 4 17 10 19
rect 4 13 5 17
rect 9 13 10 17
rect 4 -1 10 13
rect 13 5 19 19
rect 13 1 14 5
rect 18 1 19 5
rect 13 -1 19 1
rect 22 17 28 19
rect 22 13 23 17
rect 27 13 28 17
rect 22 -1 28 13
rect 31 5 37 19
rect 31 1 32 5
rect 36 1 37 5
rect 31 -1 37 1
rect 40 17 61 19
rect 40 13 41 17
rect 45 13 61 17
rect 40 -1 61 13
rect 64 6 67 19
rect 75 17 78 19
rect 77 13 78 17
rect 64 2 65 6
rect 64 -1 67 2
rect 75 -1 78 13
rect 81 10 87 19
rect 81 1 82 10
rect 86 1 87 10
rect 81 -1 87 1
rect 90 17 104 19
rect 90 13 91 17
rect 95 13 104 17
rect 90 -1 104 13
rect 107 5 113 19
rect 107 1 108 5
rect 112 1 113 5
rect 107 -1 113 1
rect 116 18 130 19
rect 116 14 117 18
rect 121 14 130 18
rect 116 -1 130 14
rect 133 5 139 19
rect 133 1 134 5
rect 138 1 139 5
rect 133 -1 139 1
rect 142 18 145 19
rect 142 14 143 18
rect 142 -1 145 14
<< ndcontact >>
rect -13 -17 -9 -13
rect 5 -24 9 -20
rect 23 -17 27 -13
rect 31 -23 35 -19
rect 47 -17 51 -13
rect 56 -23 60 -19
rect 65 -17 69 -13
rect 73 -23 77 -19
rect 91 -17 95 -13
rect 99 -23 103 -19
rect 117 -17 121 -13
rect 125 -23 129 -19
rect 143 -17 147 -13
<< pdcontact >>
rect -13 13 -9 17
rect -4 1 0 5
rect 5 13 9 17
rect 14 1 18 5
rect 23 13 27 17
rect 32 1 36 5
rect 41 13 45 17
rect 73 13 77 17
rect 65 2 69 6
rect 82 1 86 10
rect 91 13 95 17
rect 108 1 112 5
rect 117 14 121 18
rect 134 1 138 5
rect 143 14 147 18
<< polysilicon >>
rect -38 39 -36 41
rect -59 35 -57 37
rect -59 29 -57 31
rect -8 28 64 30
rect -38 25 -36 27
rect -59 21 -56 23
rect -8 19 -5 28
rect 1 19 4 20
rect 10 19 13 28
rect 19 19 22 20
rect 28 19 31 21
rect 37 19 40 21
rect 61 19 64 28
rect 78 19 81 21
rect 87 19 90 20
rect 104 19 107 21
rect 113 19 116 21
rect 130 19 133 21
rect 139 19 142 21
rect -38 12 -35 14
rect -59 -1 -56 1
rect -38 0 -35 2
rect -8 -13 -5 -1
rect 1 -13 4 -1
rect 10 -13 13 -1
rect 19 -13 22 -1
rect 28 -8 31 -1
rect 37 -2 40 -1
rect 37 -4 47 -2
rect 43 -6 47 -4
rect 28 -12 35 -8
rect 36 -13 39 -12
rect 43 -13 46 -10
rect 61 -13 64 -1
rect 78 -2 81 -1
rect 80 -6 81 -2
rect 78 -13 81 -6
rect 87 -13 90 -1
rect 104 -2 107 -1
rect 104 -13 107 -6
rect 113 -13 116 -1
rect 130 -2 133 -1
rect 131 -6 133 -2
rect 130 -13 133 -6
rect 139 -2 142 -1
rect 139 -6 141 -2
rect 139 -13 142 -6
rect -8 -25 -5 -23
rect 1 -25 4 -23
rect 10 -25 13 -23
rect 19 -25 22 -23
rect 36 -25 39 -23
rect 43 -25 46 -23
rect 61 -25 64 -23
rect 78 -25 81 -23
rect 87 -25 90 -23
rect 104 -25 107 -23
rect 113 -25 116 -23
rect 130 -25 133 -23
rect 139 -25 142 -23
<< polycontact >>
rect 0 20 4 24
rect 19 20 23 24
rect 86 20 90 24
rect 112 21 116 25
rect 35 -12 39 -8
rect 43 -10 47 -6
rect 76 -6 80 -2
rect 103 -6 107 -2
rect 127 -6 131 -2
rect 141 -6 145 -2
<< metal1 >>
rect 0 27 90 31
rect 0 24 4 27
rect 86 24 90 27
rect -9 13 5 17
rect 9 13 23 17
rect 27 13 41 17
rect 45 13 73 17
rect 77 14 91 17
rect 77 13 79 14
rect 95 14 117 17
rect 121 14 143 18
rect 100 10 145 11
rect -13 1 -4 5
rect 18 1 27 5
rect 36 1 53 5
rect -13 -2 -9 1
rect -13 -13 -9 -6
rect 23 -8 27 1
rect 23 -12 35 -8
rect 23 -13 27 -12
rect 50 -13 53 1
rect 51 -17 53 -13
rect 65 -2 69 2
rect 86 8 145 10
rect 86 7 104 8
rect 112 1 121 5
rect 65 -6 72 -2
rect 83 -3 86 1
rect 117 -2 121 1
rect 65 -13 69 -6
rect 83 -7 94 -3
rect 91 -13 94 -7
rect 117 -6 127 -2
rect 117 -13 121 -6
rect 134 -13 138 1
rect 141 -2 145 8
rect 134 -17 143 -13
rect 9 -23 31 -20
rect 35 -23 56 -20
rect 60 -23 73 -20
rect 77 -23 99 -20
rect 103 -23 125 -20
<< m2contact >>
rect 23 20 27 24
rect 108 21 112 25
rect -13 -6 -9 -2
rect 43 -6 47 -2
rect 72 -6 76 -2
rect 103 -10 107 -6
<< metal2 >>
rect 27 20 108 24
rect -9 -6 43 -2
rect 76 -6 107 -2
<< labels >>
rlabel metal1 -4 15 -4 15 1 Vdd
rlabel polycontact 2 20 3 21 1 C1?
rlabel polycontact 20 20 21 21 1 C2?
rlabel metal1 28 -22 28 -22 1 Gnd
rlabel polysilicon -7 29 -7 29 5 Iin?
<< end >>
