magic
tech scmos
timestamp 1355516091
<< nwell >>
rect 322 -274 425 -208
<< pwell >>
rect 322 -344 425 -274
<< ntransistor >>
rect 335 -295 338 -285
rect 342 -295 345 -285
rect 351 -295 354 -285
rect 358 -295 361 -285
rect 367 -295 370 -285
rect 374 -295 377 -285
rect 383 -295 386 -285
rect 390 -295 393 -285
rect 399 -291 402 -281
rect 352 -308 362 -305
rect 382 -308 392 -305
rect 402 -308 405 -298
rect 337 -333 340 -318
rect 346 -333 349 -318
rect 355 -333 358 -318
rect 364 -333 367 -318
rect 373 -333 376 -318
rect 382 -333 385 -318
rect 391 -333 394 -318
rect 400 -333 403 -318
<< ptransistor >>
rect 345 -233 365 -230
rect 384 -233 404 -230
rect 335 -264 338 -244
rect 342 -264 345 -244
rect 351 -264 354 -244
rect 358 -264 361 -244
rect 367 -264 370 -244
rect 374 -264 377 -244
rect 383 -264 386 -244
rect 390 -264 393 -244
rect 399 -268 402 -248
rect 411 -257 414 -237
<< ndiffusion >>
rect 396 -285 399 -281
rect 330 -286 335 -285
rect 334 -294 335 -286
rect 330 -295 335 -294
rect 338 -295 342 -285
rect 345 -290 351 -285
rect 345 -294 346 -290
rect 350 -294 351 -290
rect 345 -295 351 -294
rect 354 -295 358 -285
rect 361 -286 367 -285
rect 361 -294 362 -286
rect 366 -294 367 -286
rect 361 -295 367 -294
rect 370 -295 374 -285
rect 377 -290 383 -285
rect 377 -294 378 -290
rect 382 -294 383 -290
rect 377 -295 383 -294
rect 386 -295 390 -285
rect 393 -286 399 -285
rect 393 -294 394 -286
rect 398 -291 399 -286
rect 402 -282 408 -281
rect 402 -286 403 -282
rect 407 -286 408 -282
rect 402 -291 408 -286
rect 393 -295 398 -294
rect 352 -304 353 -300
rect 357 -304 362 -300
rect 352 -305 362 -304
rect 399 -299 402 -298
rect 382 -304 383 -300
rect 391 -304 392 -300
rect 382 -305 392 -304
rect 401 -307 402 -299
rect 399 -308 402 -307
rect 405 -300 409 -298
rect 405 -307 406 -300
rect 405 -308 409 -307
rect 352 -309 362 -308
rect 352 -313 353 -309
rect 361 -313 362 -309
rect 382 -309 392 -308
rect 382 -313 383 -309
rect 391 -313 392 -309
rect 332 -322 337 -318
rect 336 -326 337 -322
rect 332 -328 337 -326
rect 336 -332 337 -328
rect 332 -333 337 -332
rect 340 -319 346 -318
rect 340 -323 341 -319
rect 345 -323 346 -319
rect 340 -333 346 -323
rect 349 -326 355 -318
rect 349 -332 350 -326
rect 354 -332 355 -326
rect 349 -333 355 -332
rect 358 -319 364 -318
rect 358 -323 359 -319
rect 363 -323 364 -319
rect 358 -333 364 -323
rect 367 -319 373 -318
rect 367 -332 368 -319
rect 372 -332 373 -319
rect 367 -333 373 -332
rect 376 -319 382 -318
rect 376 -323 377 -319
rect 381 -323 382 -319
rect 376 -333 382 -323
rect 385 -326 391 -318
rect 385 -332 386 -326
rect 390 -332 391 -326
rect 385 -333 391 -332
rect 394 -319 400 -318
rect 394 -323 395 -319
rect 399 -323 400 -319
rect 394 -333 400 -323
rect 403 -322 408 -318
rect 403 -326 404 -322
rect 403 -328 408 -326
rect 403 -332 404 -328
rect 403 -333 408 -332
<< pdiffusion >>
rect 345 -229 346 -225
rect 345 -230 365 -229
rect 384 -229 385 -225
rect 384 -230 404 -229
rect 345 -234 365 -233
rect 345 -236 349 -234
rect 356 -236 365 -234
rect 384 -234 404 -233
rect 384 -236 386 -234
rect 390 -236 404 -234
rect 408 -240 411 -237
rect 410 -244 411 -240
rect 328 -245 335 -244
rect 328 -254 330 -245
rect 334 -254 335 -245
rect 328 -256 335 -254
rect 332 -264 335 -256
rect 338 -264 342 -244
rect 345 -246 351 -244
rect 345 -252 346 -246
rect 350 -252 351 -246
rect 345 -256 351 -252
rect 345 -262 346 -256
rect 350 -262 351 -256
rect 345 -264 351 -262
rect 354 -264 358 -244
rect 361 -246 367 -244
rect 361 -263 362 -246
rect 366 -263 367 -246
rect 361 -264 367 -263
rect 370 -264 374 -244
rect 377 -246 383 -244
rect 377 -252 378 -246
rect 382 -252 383 -246
rect 377 -256 383 -252
rect 377 -262 378 -256
rect 382 -262 383 -256
rect 377 -264 383 -262
rect 386 -264 390 -244
rect 393 -246 398 -244
rect 393 -262 394 -246
rect 398 -262 399 -248
rect 393 -264 399 -262
rect 396 -268 399 -264
rect 402 -261 405 -248
rect 408 -257 411 -244
rect 414 -238 417 -237
rect 414 -256 415 -238
rect 414 -257 417 -256
rect 402 -262 408 -261
rect 402 -266 403 -262
rect 407 -266 408 -262
rect 402 -268 408 -266
<< ndcontact >>
rect 330 -294 334 -286
rect 346 -294 350 -290
rect 362 -294 366 -286
rect 378 -294 382 -290
rect 394 -294 398 -286
rect 403 -286 407 -282
rect 353 -304 357 -300
rect 383 -304 391 -300
rect 397 -307 401 -299
rect 406 -307 410 -300
rect 353 -313 361 -309
rect 383 -313 391 -309
rect 332 -326 336 -322
rect 332 -332 336 -328
rect 341 -323 345 -319
rect 350 -332 354 -326
rect 359 -323 363 -319
rect 368 -332 372 -319
rect 377 -323 381 -319
rect 386 -332 390 -326
rect 395 -323 399 -319
rect 404 -326 408 -322
rect 404 -332 408 -328
<< pdcontact >>
rect 346 -229 365 -225
rect 385 -229 404 -225
rect 349 -238 356 -234
rect 386 -238 390 -234
rect 406 -244 410 -240
rect 330 -254 334 -245
rect 346 -252 350 -246
rect 346 -262 350 -256
rect 362 -263 366 -246
rect 378 -252 382 -246
rect 378 -262 382 -256
rect 394 -262 398 -246
rect 415 -256 419 -238
rect 403 -266 407 -262
<< nsubstratendiff >>
rect 416 -222 420 -218
<< psubstratepcontact >>
rect 414 -333 418 -329
<< nsubstratencontact >>
rect 412 -222 416 -218
<< polysilicon >>
rect 340 -233 345 -230
rect 365 -233 367 -230
rect 380 -233 384 -230
rect 404 -233 414 -230
rect 411 -237 414 -233
rect 335 -244 338 -242
rect 342 -244 345 -242
rect 351 -244 354 -242
rect 358 -244 361 -242
rect 367 -244 370 -242
rect 374 -244 377 -242
rect 383 -244 386 -242
rect 390 -244 393 -239
rect 399 -248 402 -246
rect 335 -272 338 -264
rect 342 -279 345 -264
rect 351 -266 354 -264
rect 358 -266 361 -264
rect 335 -285 338 -283
rect 342 -285 345 -283
rect 351 -285 354 -270
rect 367 -273 370 -264
rect 374 -266 377 -264
rect 358 -285 361 -277
rect 367 -285 370 -283
rect 374 -285 377 -270
rect 383 -279 386 -264
rect 390 -266 393 -264
rect 411 -259 414 -257
rect 399 -269 402 -268
rect 383 -285 386 -283
rect 390 -285 393 -277
rect 399 -281 402 -273
rect 399 -293 402 -291
rect 335 -297 338 -295
rect 342 -297 345 -295
rect 351 -297 354 -295
rect 358 -297 361 -295
rect 334 -301 338 -297
rect 367 -301 370 -295
rect 374 -297 377 -295
rect 383 -297 386 -295
rect 390 -297 393 -295
rect 402 -298 405 -296
rect 367 -305 368 -301
rect 346 -308 352 -305
rect 362 -308 364 -305
rect 376 -308 382 -305
rect 392 -308 396 -305
rect 393 -309 396 -308
rect 402 -309 405 -308
rect 393 -312 405 -309
rect 337 -318 340 -316
rect 346 -318 349 -316
rect 355 -318 358 -316
rect 364 -318 367 -316
rect 373 -318 376 -316
rect 382 -318 385 -316
rect 391 -318 394 -316
rect 400 -318 403 -316
rect 337 -334 340 -333
rect 346 -334 349 -333
rect 355 -334 358 -333
rect 364 -334 367 -333
rect 373 -334 376 -333
rect 382 -334 385 -333
rect 391 -334 394 -333
rect 400 -334 403 -333
rect 337 -337 403 -334
rect 337 -339 341 -337
rect 345 -339 350 -337
rect 354 -339 359 -337
rect 363 -339 377 -337
rect 381 -339 386 -337
rect 390 -339 395 -337
rect 399 -339 403 -337
<< polycontact >>
rect 340 -237 344 -233
rect 379 -237 383 -233
rect 358 -242 362 -238
rect 393 -242 397 -238
rect 334 -276 338 -272
rect 350 -270 354 -266
rect 342 -283 346 -279
rect 358 -277 362 -273
rect 366 -277 370 -273
rect 374 -270 378 -266
rect 399 -273 403 -269
rect 382 -283 386 -279
rect 390 -277 394 -273
rect 330 -301 334 -297
rect 346 -305 350 -301
rect 368 -305 372 -301
rect 376 -305 380 -301
rect 341 -341 345 -337
rect 350 -341 354 -337
rect 359 -341 363 -337
rect 377 -341 381 -337
rect 386 -341 390 -337
rect 395 -341 399 -337
<< metal1 >>
rect 322 -218 425 -211
rect 322 -222 412 -218
rect 416 -222 425 -218
rect 322 -225 425 -222
rect 322 -229 346 -225
rect 365 -229 385 -225
rect 404 -229 425 -225
rect 322 -234 334 -229
rect 330 -245 334 -234
rect 340 -246 344 -237
rect 356 -238 358 -234
rect 340 -250 346 -246
rect 324 -272 330 -262
rect 366 -251 370 -229
rect 378 -237 379 -233
rect 400 -234 425 -229
rect 378 -246 382 -237
rect 390 -242 393 -238
rect 400 -240 404 -234
rect 400 -244 406 -240
rect 400 -246 404 -244
rect 398 -251 404 -246
rect 415 -262 419 -260
rect 407 -266 411 -262
rect 354 -269 362 -266
rect 366 -269 374 -266
rect 324 -276 334 -272
rect 338 -276 358 -273
rect 324 -283 330 -276
rect 374 -276 390 -273
rect 346 -283 382 -280
rect 406 -282 411 -266
rect 415 -267 422 -262
rect 324 -311 327 -283
rect 334 -294 343 -286
rect 337 -309 343 -294
rect 330 -316 343 -309
rect 346 -301 350 -294
rect 360 -294 362 -286
rect 330 -317 337 -316
rect 322 -322 337 -317
rect 346 -319 349 -305
rect 360 -308 364 -294
rect 376 -297 382 -294
rect 407 -288 411 -282
rect 417 -285 422 -267
rect 407 -294 422 -288
rect 376 -301 380 -297
rect 394 -298 398 -294
rect 394 -299 399 -298
rect 353 -309 373 -308
rect 361 -313 373 -309
rect 367 -319 373 -313
rect 322 -326 332 -322
rect 336 -326 337 -322
rect 345 -323 359 -319
rect 367 -326 368 -319
rect 322 -328 350 -326
rect 322 -332 332 -328
rect 336 -332 350 -328
rect 354 -332 368 -326
rect 372 -326 373 -319
rect 376 -319 379 -305
rect 394 -307 397 -299
rect 394 -308 399 -307
rect 382 -309 399 -308
rect 382 -313 383 -309
rect 391 -310 399 -309
rect 391 -313 409 -310
rect 417 -311 422 -294
rect 382 -314 409 -313
rect 404 -317 409 -314
rect 376 -323 377 -319
rect 381 -323 395 -319
rect 404 -322 425 -317
rect 408 -326 425 -322
rect 372 -332 386 -326
rect 390 -328 425 -326
rect 390 -332 404 -328
rect 408 -329 425 -328
rect 408 -332 414 -329
rect 322 -333 414 -332
rect 418 -333 425 -329
rect 322 -334 425 -333
rect 322 -344 336 -334
rect 345 -341 350 -339
rect 354 -341 359 -339
rect 363 -341 377 -339
rect 381 -341 386 -339
rect 390 -341 395 -339
rect 341 -342 399 -341
rect 355 -344 359 -342
rect 381 -344 385 -342
rect 404 -344 425 -334
<< m2contact >>
rect 353 -242 358 -238
rect 346 -256 350 -252
rect 386 -242 390 -238
rect 378 -256 382 -252
rect 415 -260 419 -256
rect 362 -270 366 -266
rect 370 -277 374 -273
rect 399 -277 403 -273
rect 338 -283 342 -279
rect 330 -305 334 -301
rect 346 -290 350 -286
rect 378 -290 382 -286
rect 353 -300 357 -296
rect 368 -301 372 -297
rect 386 -300 390 -296
rect 410 -307 414 -300
<< metal2 >>
rect 338 -279 342 -207
rect 346 -286 350 -256
rect 346 -294 350 -290
rect 354 -273 358 -242
rect 362 -266 366 -207
rect 393 -242 397 -238
rect 354 -276 370 -273
rect 354 -296 358 -276
rect 378 -286 382 -256
rect 378 -294 382 -290
rect 386 -269 390 -242
rect 415 -261 419 -260
rect 410 -265 419 -261
rect 386 -272 403 -269
rect 330 -300 353 -297
rect 357 -300 358 -296
rect 386 -296 390 -272
rect 399 -273 403 -272
rect 330 -301 334 -300
rect 372 -300 386 -297
rect 410 -300 414 -265
<< labels >>
rlabel metal2 338 -208 342 -207 1 ClkB
rlabel metal2 362 -208 366 -207 1 Clk
rlabel metal1 322 -234 323 -211 1 Vpos
rlabel metal1 424 -234 425 -211 1 Vpos
rlabel metal1 322 -344 324 -317 1 Vneg
rlabel metal1 423 -344 425 -317 1 Vneg
rlabel metal1 421 -311 422 -288 1 Qb
rlabel metal1 421 -285 422 -262 1 Q
rlabel metal1 355 -344 359 -343 1 RST
rlabel metal1 324 -311 325 -262 1 D
<< end >>
