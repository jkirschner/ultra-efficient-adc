magic
tech scmos
timestamp 1355518364
<< nwell >>
rect 7 17 184 88
rect 7 9 55 17
rect 135 9 184 17
<< pwell >>
rect 55 9 134 17
rect 7 -31 184 9
<< ntransistor >>
rect 29 -9 35 3
rect 68 -5 77 3
rect 83 -5 92 3
rect 98 -5 107 3
rect 113 -5 122 3
rect 155 -9 161 3
rect 41 -24 47 -12
rect 68 -24 77 -16
rect 83 -24 92 -16
rect 98 -24 107 -16
rect 113 -24 122 -16
rect 143 -24 149 -12
<< ptransistor >>
rect 18 61 26 77
rect 32 47 92 77
rect 98 47 158 77
rect 164 61 172 77
rect 24 25 33 40
rect 39 25 48 40
rect 62 28 74 40
rect 80 28 92 40
rect 98 28 110 40
rect 116 28 128 40
rect 142 25 151 40
rect 157 25 166 40
rect 33 15 35 18
rect 155 15 157 18
<< ndiffusion >>
rect 26 1 29 3
rect 28 -8 29 1
rect 26 -9 29 -8
rect 35 1 38 3
rect 63 2 68 3
rect 35 -8 36 1
rect 67 -4 68 2
rect 63 -5 68 -4
rect 77 2 83 3
rect 77 -2 78 2
rect 82 -2 83 2
rect 77 -5 83 -2
rect 92 -2 93 3
rect 97 -2 98 3
rect 92 -5 98 -2
rect 107 2 113 3
rect 107 -2 108 2
rect 112 -2 113 2
rect 107 -5 113 -2
rect 122 2 127 3
rect 122 -4 123 2
rect 152 1 155 3
rect 122 -5 127 -4
rect 35 -9 38 -8
rect 154 -8 155 1
rect 152 -9 155 -8
rect 161 1 164 3
rect 161 -8 162 1
rect 161 -9 164 -8
rect 38 -14 41 -12
rect 40 -23 41 -14
rect 38 -24 41 -23
rect 47 -14 50 -12
rect 47 -23 48 -14
rect 140 -14 143 -12
rect 63 -17 68 -16
rect 67 -23 68 -17
rect 47 -24 50 -23
rect 63 -24 68 -23
rect 77 -19 83 -16
rect 77 -23 78 -19
rect 82 -23 83 -19
rect 77 -24 83 -23
rect 92 -24 93 -16
rect 97 -24 98 -16
rect 107 -19 113 -16
rect 107 -23 108 -19
rect 112 -23 113 -19
rect 107 -24 113 -23
rect 122 -17 127 -16
rect 122 -23 123 -17
rect 142 -23 143 -14
rect 122 -24 127 -23
rect 140 -24 143 -23
rect 149 -14 152 -12
rect 149 -23 150 -14
rect 149 -24 152 -23
<< pdiffusion >>
rect 13 75 18 77
rect 17 67 18 75
rect 13 63 18 67
rect 14 61 18 63
rect 26 76 32 77
rect 26 72 27 76
rect 31 72 32 76
rect 26 68 32 72
rect 26 61 27 68
rect 31 48 32 68
rect 29 47 32 48
rect 92 47 93 77
rect 97 47 98 77
rect 158 76 164 77
rect 158 72 159 76
rect 163 72 164 76
rect 158 68 164 72
rect 158 48 159 68
rect 163 61 164 68
rect 172 75 177 77
rect 172 67 173 75
rect 172 63 177 67
rect 172 61 176 63
rect 158 47 161 48
rect 21 38 24 40
rect 23 27 24 38
rect 21 25 24 27
rect 33 39 39 40
rect 33 35 34 39
rect 38 35 39 39
rect 33 31 39 35
rect 33 27 34 31
rect 38 27 39 31
rect 33 25 39 27
rect 48 25 49 40
rect 61 36 62 40
rect 57 32 62 36
rect 61 28 62 32
rect 74 28 75 40
rect 79 28 80 40
rect 92 28 93 40
rect 97 28 98 40
rect 110 28 111 40
rect 115 28 116 40
rect 128 36 129 40
rect 128 32 133 36
rect 128 28 129 32
rect 137 39 142 40
rect 141 26 142 39
rect 137 25 142 26
rect 151 39 157 40
rect 151 35 152 39
rect 156 35 157 39
rect 151 31 157 35
rect 151 27 152 31
rect 156 27 157 31
rect 151 25 157 27
rect 166 38 169 40
rect 166 27 167 38
rect 166 25 169 27
rect 32 15 33 18
rect 35 15 36 18
rect 154 15 155 18
rect 157 15 158 18
<< ndcontact >>
rect 24 -8 28 1
rect 36 -8 40 1
rect 63 -4 67 2
rect 78 -2 82 2
rect 93 -2 97 3
rect 108 -2 112 2
rect 123 -4 127 2
rect 150 -8 154 1
rect 162 -8 166 1
rect 36 -23 40 -14
rect 48 -23 52 -14
rect 63 -23 67 -17
rect 78 -23 82 -19
rect 93 -24 97 -16
rect 108 -23 112 -19
rect 123 -23 127 -17
rect 138 -23 142 -14
rect 150 -23 154 -14
<< pdcontact >>
rect 13 67 17 75
rect 27 72 31 76
rect 27 48 31 68
rect 93 47 97 77
rect 159 72 163 76
rect 159 48 163 68
rect 173 67 177 75
rect 19 27 23 38
rect 34 35 38 39
rect 34 27 38 31
rect 49 25 53 40
rect 57 36 61 40
rect 57 28 61 32
rect 75 28 79 40
rect 93 28 97 40
rect 111 28 115 40
rect 129 36 133 40
rect 129 28 133 32
rect 137 26 141 39
rect 152 35 156 39
rect 152 27 156 31
rect 167 27 171 38
rect 28 15 32 19
rect 36 15 40 19
rect 150 15 154 19
rect 158 15 162 19
<< psubstratepcontact >>
rect 172 -3 176 1
<< nsubstratencontact >>
rect 109 81 113 85
<< polysilicon >>
rect 18 77 26 80
rect 32 78 100 81
rect 164 79 166 80
rect 170 79 172 80
rect 104 78 158 79
rect 32 77 92 78
rect 98 77 158 78
rect 164 77 172 79
rect 18 60 26 61
rect 18 59 20 60
rect 24 59 26 60
rect 164 60 172 61
rect 164 59 166 60
rect 170 59 172 60
rect 32 45 92 47
rect 98 45 158 47
rect 24 40 33 42
rect 39 40 48 42
rect 62 40 74 42
rect 80 40 92 42
rect 98 40 110 42
rect 116 40 128 42
rect 142 40 151 42
rect 157 40 166 42
rect 62 27 74 28
rect 62 26 66 27
rect 24 23 33 25
rect 39 24 48 25
rect 39 23 43 24
rect 22 21 30 23
rect 22 8 26 21
rect 42 20 43 23
rect 47 23 48 24
rect 70 26 74 27
rect 80 26 92 28
rect 98 26 110 28
rect 116 27 128 28
rect 116 26 120 27
rect 80 23 86 26
rect 90 23 110 26
rect 124 26 128 27
rect 142 24 151 25
rect 142 23 143 24
rect 147 23 151 24
rect 157 23 166 25
rect 147 20 148 23
rect 160 21 167 23
rect 33 18 35 20
rect 33 14 35 15
rect 42 14 45 20
rect 33 11 45 14
rect 145 14 148 20
rect 155 18 157 20
rect 155 14 157 15
rect 145 11 157 14
rect 26 4 35 7
rect 29 3 35 4
rect 68 3 77 5
rect 83 4 85 5
rect 89 4 92 5
rect 83 3 92 4
rect 98 4 101 5
rect 164 8 167 21
rect 105 4 107 5
rect 98 3 107 4
rect 113 3 122 5
rect 155 3 161 7
rect 165 4 167 8
rect 68 -7 77 -5
rect 83 -7 92 -5
rect 98 -7 107 -5
rect 113 -7 122 -5
rect 29 -11 35 -9
rect 41 -11 43 -10
rect 147 -11 149 -10
rect 155 -11 161 -9
rect 41 -12 47 -11
rect 68 -15 70 -14
rect 74 -15 77 -14
rect 68 -16 77 -15
rect 83 -15 85 -14
rect 89 -15 92 -14
rect 83 -16 92 -15
rect 98 -15 101 -14
rect 105 -15 107 -14
rect 98 -16 107 -15
rect 113 -15 116 -14
rect 143 -12 149 -11
rect 120 -15 122 -14
rect 113 -16 122 -15
rect 41 -26 47 -24
rect 68 -26 77 -24
rect 83 -26 92 -24
rect 98 -26 107 -24
rect 113 -26 122 -24
rect 143 -26 149 -24
<< polycontact >>
rect 100 78 104 82
rect 166 79 170 83
rect 20 56 24 60
rect 166 56 170 60
rect 43 20 47 24
rect 66 23 70 27
rect 86 22 90 26
rect 120 23 124 27
rect 143 20 147 24
rect 22 4 26 8
rect 70 5 74 9
rect 85 4 89 8
rect 101 4 105 8
rect 116 5 120 9
rect 161 4 165 8
rect 43 -11 47 -7
rect 143 -11 147 -7
rect 70 -15 74 -11
rect 85 -15 89 -11
rect 101 -15 105 -11
rect 116 -15 120 -11
rect 144 -30 148 -26
<< metal1 >>
rect 79 82 83 88
rect 66 78 83 82
rect 41 45 45 61
rect 19 42 45 45
rect 19 38 23 42
rect 19 19 23 27
rect 43 25 49 29
rect 43 24 47 25
rect 19 15 28 19
rect 36 2 40 15
rect 50 9 53 25
rect 57 20 61 28
rect 66 31 70 78
rect 73 44 77 45
rect 73 40 79 44
rect 86 26 90 88
rect 100 82 104 88
rect 109 85 117 88
rect 113 81 117 85
rect 109 75 117 81
rect 166 83 170 88
rect 97 67 117 75
rect 118 40 122 45
rect 144 45 148 61
rect 144 42 171 45
rect 115 37 122 40
rect 93 21 97 28
rect 57 16 74 20
rect 129 20 133 28
rect 70 9 74 16
rect 116 16 133 20
rect 141 26 147 29
rect 167 38 171 42
rect 137 25 147 26
rect 89 11 101 14
rect 116 9 120 16
rect 74 5 85 8
rect 89 4 101 7
rect 105 5 116 8
rect 137 5 140 25
rect 143 24 147 25
rect 167 19 171 27
rect 162 15 171 19
rect 93 3 97 4
rect 36 1 63 2
rect 7 -8 24 1
rect 40 -2 63 1
rect 40 -4 47 -2
rect 43 -7 47 -4
rect 150 2 154 15
rect 63 -5 67 -4
rect 127 1 154 2
rect 127 -2 150 1
rect 123 -5 127 -4
rect 143 -4 150 -2
rect 7 -14 28 -8
rect 63 -8 127 -5
rect 53 -14 57 -9
rect 7 -19 36 -14
rect 7 -23 24 -19
rect 28 -23 36 -19
rect 52 -17 57 -14
rect 74 -15 85 -11
rect 89 -12 101 -11
rect 89 -15 93 -12
rect 97 -15 101 -12
rect 105 -15 116 -11
rect 133 -14 137 -9
rect 143 -7 147 -4
rect 166 -3 172 1
rect 176 -3 184 1
rect 166 -8 184 -3
rect 162 -14 184 -8
rect 52 -23 63 -17
rect 133 -17 138 -14
rect 127 -23 138 -17
rect 154 -19 184 -14
rect 154 -23 158 -19
rect 162 -23 184 -19
rect 148 -30 184 -26
<< m2contact >>
rect 13 63 17 67
rect 27 68 31 72
rect 20 52 24 56
rect 41 61 45 65
rect 34 31 38 35
rect 26 4 30 8
rect 57 32 61 36
rect 73 45 77 49
rect 66 27 70 31
rect 159 68 163 72
rect 144 61 148 65
rect 118 45 122 49
rect 173 63 177 67
rect 166 52 170 56
rect 129 32 133 36
rect 120 27 124 31
rect 93 17 97 21
rect 152 31 156 35
rect 85 11 89 15
rect 101 11 105 15
rect 50 5 54 9
rect 133 5 137 9
rect 74 -2 78 2
rect 165 4 169 8
rect 112 -2 116 2
rect 53 -9 57 -5
rect 133 -9 137 -5
rect 24 -23 28 -19
rect 93 -16 97 -12
rect 82 -22 86 -18
rect 104 -22 108 -18
rect 158 -23 162 -19
<< metal2 >>
rect 31 68 159 72
rect 13 49 16 63
rect 45 61 144 65
rect 24 52 166 56
rect 174 49 177 63
rect 13 45 73 49
rect 77 45 118 49
rect 122 45 177 49
rect 7 39 35 40
rect 57 39 133 42
rect 7 35 43 39
rect 7 31 34 35
rect 38 31 43 35
rect 57 36 61 39
rect 129 36 133 39
rect 66 33 124 36
rect 7 24 43 31
rect 66 31 70 33
rect 120 31 124 33
rect 74 24 116 30
rect 151 31 152 35
rect 156 31 184 39
rect 151 24 184 31
rect 7 19 90 24
rect 58 18 90 19
rect 100 18 184 24
rect 57 11 85 15
rect 57 9 61 11
rect 17 4 26 8
rect 54 5 61 9
rect 17 -28 21 4
rect 53 -5 57 5
rect 78 -19 82 2
rect 93 -12 97 17
rect 105 11 137 15
rect 133 9 137 11
rect 28 -22 82 -19
rect 86 -22 104 -19
rect 108 -19 112 2
rect 133 -5 137 5
rect 108 -22 158 -19
rect 28 -23 158 -22
rect 24 -25 162 -23
rect 165 -28 169 4
rect 17 -31 169 -28
<< labels >>
rlabel metal1 100 85 104 86 5 Vbias
rlabel metal1 166 85 170 86 5 Cascode
rlabel metal1 86 85 90 86 5 Vm
rlabel metal1 79 85 83 86 5 Vp
rlabel pdcontact 154 29 154 29 1 PosD
rlabel pdcontact 95 38 95 38 1 N2
rlabel metal1 95 6 95 6 1 N3
rlabel pdcontact 36 29 36 29 1 PosD
rlabel metal1 7 -23 8 1 3 Vneg
rlabel metal1 183 -23 184 1 7 Vneg
rlabel metal2 183 18 184 39 7 PosD
rlabel metal2 7 19 8 40 3 PosD
rlabel metal1 109 85 117 86 5 PosA
rlabel pdcontact 175 75 175 75 7 N1
rlabel metal2 166 -30 166 -30 1 Disable
rlabel metal1 152 8 152 8 1 Dout
rlabel metal1 183 -30 184 -26 8 Dout
<< end >>
