magic
tech scmos
timestamp 1355114294
<< nwell >>
rect 155 -297 316 -208
rect 244 -299 316 -297
<< pwell >>
rect 155 -299 244 -297
rect 155 -344 316 -299
<< ntransistor >>
rect 169 -313 172 -303
rect 178 -313 181 -303
rect 195 -313 198 -303
rect 201 -313 204 -303
rect 226 -320 229 -310
rect 233 -320 236 -310
rect 242 -320 245 -310
rect 249 -320 252 -310
rect 258 -320 261 -310
rect 265 -320 268 -310
rect 274 -320 277 -310
rect 281 -320 284 -310
rect 290 -316 293 -306
rect 174 -338 177 -328
rect 192 -338 195 -328
rect 201 -338 204 -328
rect 243 -333 253 -330
rect 273 -333 283 -330
rect 293 -333 296 -323
<< ptransistor >>
rect 174 -255 177 -235
rect 191 -255 194 -235
rect 204 -255 207 -235
rect 224 -262 227 -220
rect 233 -246 236 -220
rect 242 -246 245 -220
rect 251 -246 254 -220
rect 236 -258 256 -255
rect 263 -262 266 -220
rect 272 -246 275 -220
rect 281 -246 284 -220
rect 290 -246 293 -220
rect 275 -258 295 -255
rect 174 -289 177 -269
rect 183 -289 186 -269
rect 192 -289 195 -269
rect 201 -289 204 -269
rect 226 -289 229 -269
rect 233 -289 236 -269
rect 242 -289 245 -269
rect 249 -289 252 -269
rect 258 -289 261 -269
rect 265 -289 268 -269
rect 274 -289 277 -269
rect 281 -289 284 -269
rect 290 -293 293 -273
rect 302 -282 305 -262
<< ndiffusion >>
rect 168 -309 169 -303
rect 164 -313 169 -309
rect 172 -305 178 -303
rect 172 -313 173 -305
rect 177 -313 178 -305
rect 181 -309 182 -303
rect 181 -313 186 -309
rect 194 -309 195 -303
rect 190 -313 195 -309
rect 198 -313 201 -303
rect 204 -313 205 -303
rect 287 -310 290 -306
rect 219 -311 226 -310
rect 219 -319 221 -311
rect 225 -319 226 -311
rect 219 -320 226 -319
rect 229 -320 233 -310
rect 236 -315 242 -310
rect 236 -319 237 -315
rect 241 -319 242 -315
rect 236 -320 242 -319
rect 245 -320 249 -310
rect 252 -311 258 -310
rect 252 -319 253 -311
rect 257 -319 258 -311
rect 252 -320 258 -319
rect 261 -320 265 -310
rect 268 -315 274 -310
rect 268 -319 269 -315
rect 273 -319 274 -315
rect 268 -320 274 -319
rect 277 -320 281 -310
rect 284 -311 290 -310
rect 284 -319 285 -311
rect 289 -316 290 -311
rect 293 -307 299 -306
rect 293 -311 294 -307
rect 298 -311 299 -307
rect 293 -316 299 -311
rect 284 -320 289 -319
rect 169 -329 174 -328
rect 173 -333 174 -329
rect 169 -338 174 -333
rect 177 -329 183 -328
rect 177 -337 178 -329
rect 182 -337 183 -329
rect 177 -338 183 -337
rect 187 -329 192 -328
rect 191 -333 192 -329
rect 187 -338 192 -333
rect 195 -338 201 -328
rect 204 -329 209 -328
rect 204 -334 205 -329
rect 243 -329 244 -325
rect 248 -329 253 -325
rect 243 -330 253 -329
rect 290 -324 293 -323
rect 273 -329 274 -325
rect 282 -329 283 -325
rect 273 -330 283 -329
rect 204 -338 207 -334
rect 292 -332 293 -324
rect 290 -333 293 -332
rect 296 -325 300 -323
rect 296 -332 297 -325
rect 296 -333 300 -332
rect 243 -334 253 -333
rect 243 -338 244 -334
rect 252 -338 253 -334
rect 273 -334 283 -333
rect 273 -338 274 -334
rect 282 -338 283 -334
<< pdiffusion >>
rect 219 -227 224 -220
rect 223 -231 224 -227
rect 171 -236 174 -235
rect 173 -242 174 -236
rect 169 -246 174 -242
rect 173 -253 174 -246
rect 169 -254 174 -253
rect 171 -255 174 -254
rect 177 -236 182 -235
rect 177 -253 178 -236
rect 177 -255 182 -253
rect 186 -238 191 -235
rect 190 -242 191 -238
rect 186 -246 191 -242
rect 190 -253 191 -246
rect 186 -255 191 -253
rect 194 -241 204 -235
rect 194 -245 199 -241
rect 203 -245 204 -241
rect 194 -249 204 -245
rect 194 -253 199 -249
rect 203 -253 204 -249
rect 194 -255 204 -253
rect 207 -236 210 -235
rect 207 -253 208 -236
rect 219 -241 224 -231
rect 223 -245 224 -241
rect 207 -255 212 -253
rect 221 -262 224 -245
rect 227 -221 233 -220
rect 227 -225 228 -221
rect 232 -225 233 -221
rect 227 -234 233 -225
rect 227 -238 228 -234
rect 232 -238 233 -234
rect 227 -246 233 -238
rect 236 -227 242 -220
rect 236 -231 237 -227
rect 241 -231 242 -227
rect 236 -241 242 -231
rect 236 -245 237 -241
rect 241 -245 242 -241
rect 236 -246 242 -245
rect 245 -221 251 -220
rect 245 -225 246 -221
rect 250 -225 251 -221
rect 245 -234 251 -225
rect 245 -238 246 -234
rect 250 -238 251 -234
rect 245 -246 251 -238
rect 254 -227 263 -220
rect 254 -231 255 -227
rect 262 -231 263 -227
rect 254 -241 263 -231
rect 254 -245 255 -241
rect 262 -245 263 -241
rect 254 -246 263 -245
rect 227 -250 231 -246
rect 227 -254 228 -250
rect 236 -254 237 -250
rect 227 -262 230 -254
rect 236 -255 256 -254
rect 236 -259 256 -258
rect 236 -261 240 -259
rect 247 -261 256 -259
rect 260 -262 263 -246
rect 266 -221 272 -220
rect 266 -225 267 -221
rect 271 -225 272 -221
rect 266 -234 272 -225
rect 266 -238 267 -234
rect 271 -238 272 -234
rect 266 -246 272 -238
rect 275 -227 281 -220
rect 275 -231 276 -227
rect 280 -231 281 -227
rect 275 -241 281 -231
rect 275 -245 276 -241
rect 280 -245 281 -241
rect 275 -246 281 -245
rect 284 -221 290 -220
rect 284 -225 285 -221
rect 289 -225 290 -221
rect 284 -234 290 -225
rect 284 -238 285 -234
rect 289 -238 290 -234
rect 284 -246 290 -238
rect 293 -227 297 -220
rect 293 -231 294 -227
rect 293 -241 297 -231
rect 293 -245 294 -241
rect 293 -246 297 -245
rect 266 -250 270 -246
rect 266 -254 267 -250
rect 275 -254 276 -250
rect 266 -262 269 -254
rect 275 -255 295 -254
rect 275 -259 295 -258
rect 275 -261 277 -259
rect 281 -261 295 -259
rect 299 -265 302 -262
rect 301 -269 302 -265
rect 171 -270 174 -269
rect 173 -277 174 -270
rect 169 -281 174 -277
rect 173 -288 174 -281
rect 171 -289 174 -288
rect 177 -270 183 -269
rect 177 -288 178 -270
rect 182 -288 183 -270
rect 177 -289 183 -288
rect 186 -270 192 -269
rect 186 -277 187 -270
rect 191 -277 192 -270
rect 186 -281 192 -277
rect 186 -286 187 -281
rect 191 -286 192 -281
rect 186 -289 192 -286
rect 195 -270 201 -269
rect 195 -287 196 -270
rect 200 -287 201 -270
rect 195 -289 201 -287
rect 204 -270 207 -269
rect 219 -270 226 -269
rect 204 -288 205 -270
rect 219 -279 221 -270
rect 225 -279 226 -270
rect 204 -289 207 -288
rect 223 -289 226 -279
rect 229 -289 233 -269
rect 236 -271 242 -269
rect 236 -277 237 -271
rect 241 -277 242 -271
rect 236 -281 242 -277
rect 236 -287 237 -281
rect 241 -287 242 -281
rect 236 -289 242 -287
rect 245 -289 249 -269
rect 252 -271 258 -269
rect 252 -288 253 -271
rect 257 -288 258 -271
rect 252 -289 258 -288
rect 261 -289 265 -269
rect 268 -271 274 -269
rect 268 -277 269 -271
rect 273 -277 274 -271
rect 268 -281 274 -277
rect 268 -287 269 -281
rect 273 -287 274 -281
rect 268 -289 274 -287
rect 277 -289 281 -269
rect 284 -271 289 -269
rect 284 -287 285 -271
rect 289 -287 290 -273
rect 284 -289 290 -287
rect 287 -293 290 -289
rect 293 -286 296 -273
rect 299 -282 302 -269
rect 305 -263 308 -262
rect 305 -281 306 -263
rect 305 -282 308 -281
rect 293 -287 299 -286
rect 293 -291 294 -287
rect 298 -291 299 -287
rect 293 -293 299 -291
<< ndcontact >>
rect 164 -309 168 -303
rect 173 -313 177 -305
rect 182 -309 186 -303
rect 190 -309 194 -303
rect 205 -313 209 -303
rect 221 -319 225 -311
rect 237 -319 241 -315
rect 253 -319 257 -311
rect 269 -319 273 -315
rect 285 -319 289 -311
rect 294 -311 298 -307
rect 169 -333 173 -329
rect 178 -337 182 -329
rect 187 -333 191 -329
rect 205 -334 209 -329
rect 244 -329 248 -325
rect 274 -329 282 -325
rect 288 -332 292 -324
rect 297 -332 301 -325
rect 244 -338 252 -334
rect 274 -338 282 -334
<< pdcontact >>
rect 219 -231 223 -227
rect 169 -242 173 -236
rect 169 -253 173 -246
rect 178 -253 182 -236
rect 186 -242 190 -238
rect 186 -253 190 -246
rect 199 -245 203 -241
rect 199 -253 203 -249
rect 208 -253 212 -236
rect 219 -245 223 -241
rect 228 -225 232 -221
rect 228 -238 232 -234
rect 237 -231 241 -227
rect 237 -245 241 -241
rect 246 -225 250 -221
rect 246 -238 250 -234
rect 255 -231 262 -227
rect 255 -245 262 -241
rect 228 -254 232 -250
rect 237 -254 256 -250
rect 240 -263 247 -259
rect 267 -225 271 -221
rect 267 -238 271 -234
rect 276 -231 280 -227
rect 276 -245 280 -241
rect 285 -225 289 -221
rect 285 -238 289 -234
rect 294 -231 298 -227
rect 294 -245 298 -241
rect 267 -254 271 -250
rect 276 -254 295 -250
rect 277 -263 281 -259
rect 297 -269 301 -265
rect 169 -277 173 -270
rect 169 -288 173 -281
rect 178 -288 182 -270
rect 187 -277 191 -270
rect 187 -286 191 -281
rect 196 -287 200 -270
rect 205 -288 209 -270
rect 221 -279 225 -270
rect 237 -277 241 -271
rect 237 -287 241 -281
rect 253 -288 257 -271
rect 269 -277 273 -271
rect 269 -287 273 -281
rect 285 -287 289 -271
rect 306 -281 310 -263
rect 294 -291 298 -287
<< psubstratepdiff >>
rect 222 -336 226 -332
<< nsubstratendiff >>
rect 307 -221 311 -217
<< psubstratepcontact >>
rect 226 -336 230 -332
<< nsubstratencontact >>
rect 303 -221 307 -217
<< polysilicon >>
rect 224 -218 228 -216
rect 232 -218 237 -216
rect 241 -218 246 -216
rect 250 -218 267 -216
rect 271 -218 276 -216
rect 280 -218 285 -216
rect 289 -218 293 -216
rect 224 -219 293 -218
rect 224 -220 227 -219
rect 233 -220 236 -219
rect 242 -220 245 -219
rect 251 -220 254 -219
rect 263 -220 266 -219
rect 272 -220 275 -219
rect 281 -220 284 -219
rect 290 -220 293 -219
rect 174 -235 177 -233
rect 191 -235 194 -233
rect 204 -235 207 -233
rect 174 -269 177 -255
rect 191 -256 194 -255
rect 204 -256 207 -255
rect 181 -259 194 -256
rect 206 -260 207 -256
rect 233 -248 236 -246
rect 242 -248 245 -246
rect 251 -248 254 -246
rect 231 -258 236 -255
rect 256 -258 258 -255
rect 194 -267 195 -263
rect 224 -264 227 -262
rect 272 -248 275 -246
rect 281 -248 284 -246
rect 290 -248 293 -246
rect 270 -258 275 -255
rect 295 -258 305 -255
rect 263 -264 266 -262
rect 302 -262 305 -258
rect 183 -269 186 -267
rect 192 -269 195 -267
rect 201 -269 204 -267
rect 226 -269 229 -267
rect 233 -269 236 -267
rect 242 -269 245 -267
rect 249 -269 252 -267
rect 258 -269 261 -267
rect 265 -269 268 -267
rect 274 -269 277 -267
rect 281 -269 284 -264
rect 290 -273 293 -271
rect 174 -291 177 -289
rect 168 -294 177 -291
rect 183 -291 186 -289
rect 168 -295 172 -294
rect 169 -303 172 -295
rect 183 -295 184 -291
rect 183 -297 186 -295
rect 178 -300 186 -297
rect 192 -298 195 -289
rect 178 -303 181 -300
rect 192 -301 198 -298
rect 195 -303 198 -301
rect 201 -303 204 -289
rect 226 -297 229 -289
rect 233 -304 236 -289
rect 242 -291 245 -289
rect 249 -291 252 -289
rect 226 -310 229 -308
rect 233 -310 236 -308
rect 242 -310 245 -295
rect 258 -298 261 -289
rect 265 -291 268 -289
rect 249 -310 252 -302
rect 258 -310 261 -308
rect 265 -310 268 -295
rect 274 -304 277 -289
rect 281 -291 284 -289
rect 302 -284 305 -282
rect 290 -294 293 -293
rect 274 -310 277 -308
rect 281 -310 284 -302
rect 290 -306 293 -298
rect 169 -324 172 -313
rect 178 -315 181 -313
rect 195 -316 198 -313
rect 201 -315 204 -313
rect 197 -320 198 -316
rect 290 -318 293 -316
rect 226 -322 229 -320
rect 233 -322 236 -320
rect 242 -322 245 -320
rect 249 -322 252 -320
rect 185 -324 189 -322
rect 169 -327 177 -324
rect 185 -327 195 -324
rect 202 -326 203 -322
rect 174 -328 177 -327
rect 192 -328 195 -327
rect 201 -327 207 -326
rect 201 -328 204 -327
rect 258 -326 261 -320
rect 265 -322 268 -320
rect 274 -322 277 -320
rect 281 -322 284 -320
rect 293 -323 296 -321
rect 258 -330 259 -326
rect 237 -333 243 -330
rect 253 -333 255 -330
rect 267 -333 273 -330
rect 283 -333 287 -330
rect 284 -334 287 -333
rect 293 -334 296 -333
rect 284 -337 296 -334
rect 174 -340 177 -338
rect 192 -340 195 -338
rect 201 -340 204 -338
<< polycontact >>
rect 228 -218 232 -214
rect 237 -218 241 -214
rect 246 -218 250 -214
rect 267 -218 271 -214
rect 276 -218 280 -214
rect 285 -218 289 -214
rect 181 -263 185 -259
rect 202 -260 206 -256
rect 231 -262 235 -258
rect 190 -267 194 -263
rect 270 -262 274 -258
rect 249 -267 253 -263
rect 284 -267 288 -263
rect 164 -295 168 -291
rect 184 -295 188 -291
rect 204 -299 208 -295
rect 225 -301 229 -297
rect 241 -295 245 -291
rect 233 -308 237 -304
rect 249 -302 253 -298
rect 257 -302 261 -298
rect 265 -295 269 -291
rect 290 -298 294 -294
rect 273 -308 277 -304
rect 281 -302 285 -298
rect 185 -322 189 -318
rect 193 -320 197 -316
rect 203 -326 207 -322
rect 225 -326 229 -322
rect 237 -330 241 -326
rect 259 -330 263 -326
rect 267 -330 271 -326
<< metal1 >>
rect 155 -234 160 -211
rect 218 -227 223 -211
rect 242 -213 246 -208
rect 228 -214 289 -213
rect 232 -216 237 -214
rect 241 -216 246 -214
rect 250 -216 267 -214
rect 271 -216 276 -214
rect 280 -216 285 -214
rect 294 -216 316 -211
rect 293 -217 316 -216
rect 293 -221 303 -217
rect 307 -221 316 -217
rect 232 -224 246 -221
rect 254 -227 263 -221
rect 271 -224 285 -221
rect 293 -227 316 -221
rect 218 -231 219 -227
rect 223 -231 237 -228
rect 254 -228 255 -227
rect 241 -231 255 -228
rect 262 -228 263 -227
rect 262 -231 276 -228
rect 293 -228 294 -227
rect 280 -231 294 -228
rect 298 -231 316 -227
rect 218 -232 224 -231
rect 179 -235 196 -232
rect 179 -236 182 -235
rect 193 -256 196 -235
rect 217 -241 224 -232
rect 232 -238 246 -234
rect 254 -241 263 -231
rect 293 -234 316 -231
rect 271 -238 285 -234
rect 293 -241 307 -234
rect 217 -244 219 -241
rect 212 -245 219 -244
rect 223 -245 237 -241
rect 241 -245 255 -241
rect 262 -245 276 -241
rect 280 -245 294 -241
rect 298 -245 307 -241
rect 212 -247 307 -245
rect 212 -253 225 -247
rect 236 -250 264 -247
rect 275 -250 307 -247
rect 191 -259 196 -256
rect 178 -263 181 -259
rect 191 -263 194 -259
rect 157 -291 161 -264
rect 178 -270 182 -263
rect 199 -263 206 -260
rect 199 -270 202 -263
rect 221 -270 225 -253
rect 200 -274 202 -270
rect 157 -295 164 -291
rect 157 -313 161 -295
rect 178 -298 181 -288
rect 178 -301 186 -298
rect 182 -303 186 -301
rect 197 -303 200 -287
rect 209 -279 221 -270
rect 236 -254 237 -250
rect 256 -254 264 -250
rect 275 -254 276 -250
rect 295 -254 307 -250
rect 228 -258 232 -254
rect 228 -262 231 -258
rect 228 -271 232 -262
rect 247 -263 249 -259
rect 228 -275 237 -271
rect 216 -297 220 -286
rect 257 -276 261 -254
rect 267 -258 271 -254
rect 267 -262 270 -258
rect 267 -271 272 -262
rect 281 -267 284 -263
rect 291 -265 295 -254
rect 306 -263 313 -262
rect 291 -269 297 -265
rect 291 -271 295 -269
rect 267 -273 269 -271
rect 289 -276 295 -271
rect 310 -285 313 -263
rect 298 -288 300 -287
rect 298 -291 313 -288
rect 245 -294 253 -291
rect 257 -294 265 -291
rect 216 -302 225 -297
rect 229 -301 249 -298
rect 265 -301 281 -298
rect 164 -317 168 -313
rect 155 -321 168 -317
rect 183 -318 186 -309
rect 197 -307 205 -303
rect 203 -313 205 -307
rect 212 -307 225 -302
rect 155 -329 173 -321
rect 183 -322 185 -318
rect 197 -320 198 -316
rect 155 -344 169 -329
rect 195 -337 198 -320
rect 203 -322 207 -313
rect 212 -316 216 -307
rect 237 -308 273 -305
rect 297 -307 313 -291
rect 298 -311 308 -307
rect 312 -311 313 -307
rect 210 -319 216 -316
rect 219 -319 221 -311
rect 210 -329 213 -319
rect 219 -322 222 -319
rect 209 -334 213 -329
rect 217 -329 222 -322
rect 237 -326 241 -319
rect 251 -319 253 -311
rect 217 -332 234 -329
rect 217 -336 226 -332
rect 230 -333 234 -332
rect 251 -333 255 -319
rect 267 -322 273 -319
rect 267 -326 271 -322
rect 285 -323 289 -319
rect 285 -324 290 -323
rect 285 -332 288 -324
rect 301 -332 305 -329
rect 285 -333 290 -332
rect 230 -334 290 -333
rect 230 -336 244 -334
rect 217 -337 244 -336
rect 178 -340 198 -337
rect 213 -338 244 -337
rect 252 -338 274 -334
rect 282 -335 290 -334
rect 308 -335 316 -317
rect 282 -338 316 -335
rect 213 -344 316 -338
<< m2contact >>
rect 160 -234 164 -211
rect 213 -232 218 -211
rect 169 -246 173 -242
rect 186 -246 190 -242
rect 199 -241 203 -237
rect 199 -249 203 -245
rect 169 -281 173 -277
rect 187 -281 191 -277
rect 188 -295 192 -291
rect 244 -267 249 -263
rect 237 -281 241 -277
rect 216 -286 220 -282
rect 208 -299 212 -295
rect 277 -267 281 -263
rect 269 -281 273 -277
rect 306 -285 310 -281
rect 253 -295 257 -291
rect 261 -302 265 -298
rect 290 -302 294 -298
rect 164 -313 168 -309
rect 190 -313 194 -309
rect 187 -329 191 -325
rect 169 -344 173 -333
rect 229 -308 233 -304
rect 308 -311 312 -307
rect 237 -315 241 -311
rect 229 -326 233 -322
rect 269 -315 273 -311
rect 244 -325 248 -321
rect 259 -326 263 -322
rect 277 -325 281 -321
rect 301 -329 305 -325
rect 209 -344 213 -337
<< metal2 >>
rect 164 -232 213 -211
rect 164 -234 191 -232
rect 169 -242 191 -234
rect 173 -246 186 -242
rect 190 -246 191 -242
rect 169 -277 191 -246
rect 199 -244 203 -241
rect 199 -245 220 -244
rect 203 -249 220 -245
rect 173 -281 187 -277
rect 216 -282 220 -249
rect 188 -291 226 -289
rect 192 -292 226 -291
rect 168 -313 190 -309
rect 164 -325 194 -313
rect 164 -329 187 -325
rect 191 -329 194 -325
rect 164 -333 194 -329
rect 164 -344 169 -333
rect 173 -337 194 -333
rect 208 -331 212 -299
rect 222 -329 226 -292
rect 229 -304 233 -208
rect 237 -311 241 -281
rect 237 -319 241 -315
rect 245 -298 249 -267
rect 253 -291 257 -208
rect 284 -267 288 -263
rect 245 -301 261 -298
rect 245 -321 249 -301
rect 269 -311 273 -281
rect 269 -319 273 -315
rect 277 -294 281 -267
rect 301 -285 306 -281
rect 277 -297 294 -294
rect 233 -325 244 -322
rect 248 -325 249 -321
rect 277 -321 281 -297
rect 290 -298 294 -297
rect 263 -325 277 -322
rect 301 -325 305 -285
rect 208 -334 219 -331
rect 222 -333 305 -329
rect 216 -337 219 -334
rect 308 -337 312 -311
rect 173 -344 209 -337
rect 216 -340 312 -337
rect 216 -341 311 -340
<< labels >>
rlabel metal1 314 -344 316 -317 1 Vneg
rlabel metal1 315 -234 316 -211 1 Vpos
rlabel metal1 312 -311 313 -288 1 Qb
rlabel metal2 229 -209 233 -208 1 ClkB
rlabel metal2 253 -209 257 -208 1 Clk
rlabel metal1 242 -209 246 -208 1 RstB
rlabel pwell 212 -344 214 -317 3 Vneg
rlabel metal1 312 -285 313 -262 1 Q
rlabel metal1 157 -313 158 -264 3 T
rlabel metal1 155 -344 156 -317 3 Vneg
rlabel metal1 155 -234 156 -211 3 Vpos
<< end >>
