magic
tech scmos
timestamp 1355540337
<< nwell >>
rect -8 27 11 68
rect -8 -8 4 27
rect -8 -22 11 -8
rect -1 -41 11 -22
rect -1 -60 55 -41
rect 9 -63 55 -60
rect 154 -4 169 64
rect 268 -44 283 22
rect 386 -32 397 22
rect 383 -55 399 -32
rect 500 -40 585 19
rect 500 -55 523 -40
rect 577 -41 585 -40
rect 386 -69 397 -55
rect 688 -69 697 22
rect 800 20 808 22
rect 800 -33 806 20
rect 909 -15 924 19
rect 908 -32 990 -15
rect 797 -55 808 -33
rect 908 -42 989 -32
rect 905 -46 989 -42
rect 908 -47 989 -46
rect 970 -49 989 -47
rect 1037 -46 1043 19
rect 1145 -4 1191 20
rect 1037 -50 1045 -46
rect 800 -69 806 -55
rect 1175 -155 1191 -4
rect 1170 -156 1191 -155
rect 1160 -174 1191 -156
rect 1161 -180 1191 -174
rect 154 -331 185 -228
rect 259 -276 276 -275
rect 311 -290 343 -275
rect 153 -395 185 -331
rect 299 -338 343 -290
rect 304 -386 343 -338
rect 272 -395 343 -386
rect 392 -395 425 -277
rect 470 -395 501 -277
rect 542 -395 578 -277
rect 622 -395 654 -277
rect 727 -395 759 -276
rect 797 -387 826 -333
rect 89 -397 759 -395
rect 797 -397 829 -387
rect 875 -397 906 -276
rect 1175 -227 1191 -180
rect 960 -397 992 -277
rect 1161 -396 1193 -291
rect 1128 -397 1196 -396
rect 89 -422 1196 -397
<< pwell >>
rect 139 -44 154 0
rect 139 -83 165 -44
rect 86 -101 165 -83
rect 86 -113 177 -101
rect 268 -113 283 -69
rect 386 -113 397 -69
rect 500 -71 523 -56
rect 571 -71 585 -69
rect 500 -113 585 -71
rect 688 -113 697 -69
rect 800 -113 806 -69
rect 909 -79 922 -65
rect 970 -79 989 -50
rect 1036 -79 1043 -53
rect 909 -113 1043 -79
rect 1135 -113 1146 -112
rect 86 -114 1146 -113
rect 134 -120 1146 -114
rect 121 -155 1146 -120
rect 121 -179 1160 -155
rect 121 -180 1145 -179
rect 121 -204 1148 -180
rect 121 -245 153 -204
rect 133 -276 153 -245
rect 212 -276 244 -204
rect 279 -276 311 -204
rect 212 -290 255 -276
rect 360 -277 392 -204
rect 438 -232 468 -204
rect 438 -246 457 -232
rect 511 -277 542 -204
rect 590 -277 622 -204
rect 695 -277 727 -204
rect 240 -386 272 -338
rect 762 -285 794 -204
rect 843 -276 875 -204
rect 762 -331 793 -285
rect 765 -332 781 -331
rect 765 -387 793 -332
rect 928 -277 960 -204
rect 1129 -396 1161 -291
<< ntransistor >>
rect 1145 -316 1155 -313
<< ptransistor >>
rect 1167 -316 1187 -313
<< ndiffusion >>
rect 1149 -312 1155 -310
rect 1145 -313 1155 -312
rect 1145 -317 1155 -316
rect 1145 -319 1151 -317
<< pdiffusion >>
rect 1167 -311 1176 -310
rect 1186 -311 1187 -310
rect 1167 -313 1187 -311
rect 1167 -317 1187 -316
rect 1167 -319 1168 -317
rect 1172 -319 1187 -317
<< ndcontact >>
rect 1145 -312 1149 -308
rect 1151 -321 1155 -317
<< pdcontact >>
rect 1176 -311 1186 -307
rect 1168 -321 1172 -317
<< psubstratepcontact >>
rect 1134 -326 1138 -322
<< nsubstratencontact >>
rect 1185 -331 1189 -327
<< polysilicon >>
rect 1143 -316 1145 -313
rect 1155 -314 1158 -313
rect 1162 -314 1167 -313
rect 1155 -316 1167 -314
rect 1187 -316 1189 -313
<< polycontact >>
rect 1158 -314 1162 -310
<< metal1 >>
rect -8 57 11 68
rect -8 -8 4 57
rect 73 55 81 62
rect 154 46 165 64
rect 519 52 977 56
rect 11 0 79 2
rect -8 -22 11 -8
rect -1 -41 11 -22
rect -1 -60 55 -41
rect 9 -63 55 -60
rect -10 -84 55 -80
rect 141 -87 154 0
rect 161 -4 165 46
rect 172 26 176 43
rect 181 26 185 36
rect 205 26 209 29
rect 299 26 303 36
rect 312 26 316 45
rect 413 26 417 36
rect 426 22 430 45
rect 519 26 523 52
rect 601 26 605 36
rect 614 22 618 45
rect 713 26 717 36
rect 726 22 730 45
rect 822 26 826 36
rect 835 22 839 45
rect 268 -4 283 19
rect 386 -4 397 19
rect 500 -4 585 19
rect 688 -4 697 19
rect 800 -4 806 19
rect 909 -4 924 19
rect 265 -55 285 -32
rect 383 -55 399 -32
rect 512 -40 571 -4
rect 913 -32 924 -4
rect 973 -3 977 52
rect 1059 26 1063 36
rect 1072 22 1076 45
rect 970 -32 990 -15
rect 1037 -25 1043 19
rect 1145 -4 1191 20
rect 1037 -29 1042 -25
rect 1150 -31 1156 -15
rect 554 -57 587 -53
rect 685 -55 699 -32
rect 797 -55 808 -33
rect 905 -46 922 -42
rect 973 -45 977 -40
rect 970 -49 977 -45
rect 1023 -53 1045 -42
rect 1143 -55 1156 -31
rect 519 -58 523 -57
rect 265 -63 279 -58
rect 265 -75 272 -63
rect 278 -75 279 -63
rect 265 -81 279 -75
rect 383 -62 394 -58
rect 383 -74 388 -62
rect 393 -74 394 -62
rect 497 -65 523 -58
rect 685 -60 694 -58
rect 383 -81 394 -74
rect 141 -101 165 -87
rect 103 -114 177 -101
rect 141 -120 165 -114
rect 268 -114 283 -87
rect 386 -114 397 -87
rect 500 -88 571 -71
rect 685 -79 687 -60
rect 692 -79 694 -60
rect 685 -81 694 -79
rect 909 -79 922 -65
rect 970 -79 989 -64
rect 909 -87 1037 -79
rect 500 -114 585 -88
rect 688 -114 697 -87
rect 800 -114 806 -87
rect 909 -114 1043 -87
rect 372 -120 1145 -114
rect 121 -134 1145 -120
rect 121 -141 385 -134
rect 121 -245 140 -141
rect 150 -228 154 -158
rect 212 -259 228 -141
rect 238 -231 242 -158
rect 245 -228 249 -208
rect 279 -259 295 -141
rect 305 -228 309 -219
rect 312 -228 316 -196
rect 360 -246 379 -141
rect 388 -204 393 -153
rect 389 -231 393 -208
rect 438 -246 457 -134
rect 467 -248 471 -166
rect 511 -236 524 -134
rect 534 -229 538 -208
rect 541 -229 545 -180
rect 548 -229 552 -219
rect 590 -260 606 -134
rect 616 -229 620 -166
rect 623 -229 627 -173
rect 687 -215 692 -144
rect 695 -260 711 -134
rect 721 -229 725 -166
rect 728 -229 732 -180
rect 149 -388 153 -276
rect 167 -400 185 -276
rect 212 -285 228 -276
rect 259 -281 276 -275
rect 326 -281 343 -275
rect 271 -284 343 -281
rect 212 -290 255 -285
rect 290 -290 304 -284
rect 389 -386 393 -277
rect 89 -401 255 -400
rect 286 -401 304 -386
rect 406 -400 425 -277
rect 467 -382 471 -277
rect 484 -400 501 -277
rect 541 -384 545 -277
rect 562 -400 574 -277
rect 620 -382 624 -276
rect 637 -400 654 -277
rect 742 -400 759 -276
rect 762 -300 780 -134
rect 792 -169 797 -145
rect 828 -260 833 -173
rect 869 -228 873 -173
rect 876 -228 880 -180
rect 928 -246 946 -134
rect 980 -176 985 -143
rect 1130 -180 1145 -134
rect 1175 -179 1191 -4
rect 1158 -180 1162 -179
rect 957 -229 961 -180
rect 765 -340 781 -330
rect 791 -339 795 -333
rect 873 -374 877 -276
rect 812 -400 829 -387
rect 890 -400 906 -276
rect 957 -382 961 -277
rect 974 -400 992 -277
rect 1129 -308 1148 -291
rect 1129 -312 1145 -308
rect 1158 -310 1162 -291
rect 1129 -322 1148 -312
rect 1175 -307 1193 -291
rect 1175 -311 1176 -307
rect 1186 -311 1193 -307
rect 1155 -321 1168 -317
rect 1129 -326 1134 -322
rect 1138 -326 1148 -322
rect 1129 -396 1148 -326
rect 1158 -335 1162 -321
rect 1175 -327 1193 -311
rect 1175 -331 1185 -327
rect 1189 -331 1193 -327
rect 1175 -397 1193 -331
rect 1175 -400 1196 -397
rect 355 -401 1196 -400
rect 89 -422 1196 -401
<< m2contact >>
rect 114 29 118 33
rect 154 29 158 33
rect 8 25 12 29
rect 103 -77 107 -73
rect -14 -84 -10 -80
rect 103 -84 107 -80
rect 172 43 176 47
rect 312 45 316 49
rect 172 22 176 26
rect 181 36 185 40
rect 299 36 303 40
rect 181 22 185 26
rect 205 29 209 33
rect 205 22 209 26
rect 299 22 303 26
rect 426 45 430 49
rect 312 22 316 26
rect 413 36 417 40
rect 413 22 417 26
rect 614 45 618 49
rect 519 22 523 26
rect 601 36 605 40
rect 601 22 605 26
rect 726 45 730 49
rect 713 36 717 40
rect 713 22 717 26
rect 835 45 839 49
rect 822 36 826 40
rect 822 22 826 26
rect 164 -60 168 -34
rect 1072 45 1076 49
rect 1059 36 1063 40
rect 1059 22 1063 26
rect 973 -7 977 -3
rect 1150 -15 1156 -11
rect 519 -54 523 -50
rect 973 -40 977 -36
rect 985 -47 989 -43
rect 918 -53 922 -49
rect 985 -54 989 -50
rect 272 -75 278 -63
rect 388 -74 393 -62
rect 492 -78 496 -66
rect 103 -91 107 -87
rect 198 -117 202 -113
rect 687 -79 692 -60
rect 792 -78 797 -59
rect 906 -62 910 -58
rect 1138 -79 1142 -60
rect 150 -158 154 -154
rect 238 -158 242 -154
rect 245 -208 249 -204
rect 312 -196 316 -192
rect 305 -219 309 -215
rect 388 -153 393 -146
rect 388 -208 393 -204
rect 467 -166 471 -162
rect 541 -180 545 -176
rect 534 -208 538 -204
rect 548 -219 552 -215
rect 687 -144 692 -140
rect 616 -166 620 -162
rect 623 -173 627 -169
rect 687 -219 692 -215
rect 721 -166 725 -162
rect 728 -180 732 -176
rect 242 -276 246 -272
rect 149 -392 153 -388
rect 309 -276 313 -272
rect 265 -294 269 -290
rect 272 -294 276 -290
rect 269 -390 273 -386
rect 389 -390 393 -386
rect 467 -386 471 -382
rect 541 -388 545 -384
rect 620 -386 624 -382
rect 725 -281 729 -277
rect 792 -145 797 -141
rect 792 -173 797 -169
rect 828 -173 833 -169
rect 869 -173 873 -169
rect 876 -180 880 -176
rect 980 -143 985 -139
rect 957 -180 961 -176
rect 980 -180 985 -176
rect 1158 -179 1162 -175
rect 828 -264 833 -260
rect 791 -285 795 -281
rect 798 -339 802 -335
rect 873 -378 877 -374
rect 795 -391 799 -387
rect 957 -386 961 -382
rect 1158 -396 1162 -335
<< metal2 >>
rect 466 59 1156 63
rect 466 56 473 59
rect 290 52 473 56
rect 290 47 295 52
rect 176 43 295 47
rect 316 45 426 49
rect 430 45 614 49
rect 618 45 726 49
rect 730 45 835 49
rect 839 45 1072 49
rect 1076 45 1091 49
rect 114 36 181 40
rect 185 36 299 40
rect 303 36 413 40
rect 417 36 601 40
rect 605 36 713 40
rect 717 36 822 40
rect 826 36 1059 40
rect 1063 36 1103 40
rect 114 33 118 36
rect 158 29 205 33
rect 209 29 1099 33
rect -14 25 8 29
rect -14 -80 -10 25
rect 164 22 172 26
rect 323 22 327 29
rect 437 22 441 29
rect 625 22 629 29
rect 737 22 741 29
rect 846 22 850 29
rect 1083 22 1087 29
rect 164 -34 168 22
rect 519 -50 523 22
rect 973 -36 977 -7
rect 1150 -11 1156 59
rect 918 -47 985 -43
rect 918 -49 922 -47
rect 971 -54 985 -50
rect 971 -58 975 -54
rect 107 -77 130 -73
rect 107 -84 122 -80
rect 107 -91 115 -87
rect 111 -176 115 -91
rect 118 -169 122 -84
rect 126 -162 130 -77
rect 272 -154 278 -75
rect 388 -146 393 -74
rect 492 -121 496 -78
rect 141 -158 150 -154
rect 154 -158 238 -154
rect 242 -158 280 -154
rect 492 -162 497 -121
rect 687 -140 692 -79
rect 792 -141 797 -78
rect 910 -62 975 -58
rect 906 -117 910 -62
rect 980 -139 985 -54
rect 1138 -107 1142 -79
rect 1138 -111 1162 -107
rect 126 -166 467 -162
rect 471 -166 616 -162
rect 620 -166 721 -162
rect 725 -166 1069 -162
rect 118 -173 623 -169
rect 627 -173 792 -169
rect 797 -173 828 -169
rect 833 -173 869 -169
rect 873 -173 1069 -169
rect 1158 -170 1162 -111
rect 1125 -171 1162 -170
rect 1085 -175 1162 -171
rect 111 -180 541 -176
rect 545 -180 728 -176
rect 732 -180 876 -176
rect 880 -180 957 -176
rect 961 -180 980 -176
rect 985 -180 1069 -176
rect 1085 -179 1158 -175
rect 1085 -192 1098 -179
rect 141 -196 312 -192
rect 316 -196 1098 -192
rect 141 -208 245 -204
rect 249 -208 388 -204
rect 393 -208 534 -204
rect 538 -208 1069 -204
rect 141 -219 305 -215
rect 309 -219 548 -215
rect 552 -219 687 -215
rect 692 -219 1069 -215
rect 242 -281 246 -276
rect 309 -278 313 -276
rect 272 -281 313 -278
rect 729 -281 794 -280
rect 242 -285 269 -281
rect 265 -290 269 -285
rect 272 -284 279 -281
rect 272 -290 276 -284
rect 725 -285 791 -281
rect 149 -431 153 -392
rect 269 -427 273 -390
rect 389 -439 393 -390
rect 467 -441 471 -386
rect 541 -436 545 -388
rect 620 -432 624 -386
rect 725 -431 729 -285
rect 828 -335 833 -264
rect 802 -339 833 -335
rect 873 -374 877 -373
rect 795 -431 799 -391
rect 873 -429 877 -378
rect 957 -428 961 -386
rect 1158 -432 1162 -396
use SPDT  SPDT_0
timestamp 1355531441
transform 1 0 -27 0 1 0
box 38 1 105 68
use NOT  NOT_0
timestamp 1355475633
transform 1 0 83 0 1 23
box -5 -23 43 41
use NOT  NOT_1
timestamp 1355475633
transform 1 0 111 0 1 23
box -5 -23 43 41
use NAND3  NAND3_0
timestamp 1355475992
transform -1 0 91 0 1 -72
box -12 -42 36 26
use ResetFlipFlop_High_Layout  ResetFlipFlop_High_Layout_0
timestamp 1355516091
transform 1 0 -157 0 1 230
box 322 -344 425 -207
use ResetFlipFlop_Low_Layout  ResetFlipFlop_Low_Layout_0
timestamp 1354992098
transform 1 0 70 0 1 230
box 213 -344 316 -208
use ResetFlipFlop_Low_Layout  ResetFlipFlop_Low_Layout_1
timestamp 1354992098
transform 1 0 184 0 1 230
box 213 -344 316 -208
use NAND  NAND_0
timestamp 1355475793
transform 1 0 539 0 1 -85
box -16 -2 32 62
use ResetFlipFlop_Low_Layout  ResetFlipFlop_Low_Layout_2
timestamp 1354992098
transform 1 0 372 0 1 230
box 213 -344 316 -208
use ResetFlipFlop_Low_Layout  ResetFlipFlop_Low_Layout_3
timestamp 1354992098
transform 1 0 484 0 1 230
box 213 -344 316 -208
use ResetFlipFlop_Low_Layout  ResetFlipFlop_Low_Layout_4
timestamp 1354992098
transform 1 0 593 0 1 230
box 213 -344 316 -208
use NAND  NAND_1
timestamp 1355475793
transform 1 0 938 0 1 -77
box -16 -2 32 62
use NOR  NOR_0
timestamp 1355475848
transform 1 0 1003 0 1 -57
box -14 -22 34 42
use ResetFlipFlop_Low_Layout  ResetFlipFlop_Low_Layout_5
timestamp 1354992098
transform 1 0 830 0 1 230
box 213 -344 316 -208
use NOT  NOT_2
timestamp 1355475633
transform 0 1 1152 -1 0 -184
box -5 -23 43 41
use NOT  NOT_6
timestamp 1355475633
transform 0 1 144 -1 0 -233
box -5 -23 43 41
use NAND  NAND_2
timestamp 1355475793
transform 0 1 214 -1 0 -244
box -16 -2 32 62
use NAND  NAND_3
timestamp 1355475793
transform 0 1 281 -1 0 -244
box -16 -2 32 62
use NOT  NOT_8
timestamp 1355475633
transform 0 1 383 -1 0 -234
box -5 -23 43 41
use NOT  NOT_9
timestamp 1355475633
transform 0 1 461 -1 0 -234
box -5 -23 43 41
use NAND3  NAND3_1
timestamp 1355475992
transform 0 1 553 -1 0 -241
box -12 -42 36 26
use NAND  NAND_4
timestamp 1355475793
transform 0 1 592 -1 0 -245
box -16 -2 32 62
use NAND  NAND_5
timestamp 1355475793
transform 0 1 697 -1 0 -245
box -16 -2 32 62
use NAND  NAND_7
timestamp 1355475793
transform 0 1 845 -1 0 -244
box -16 -2 32 62
use NOT  NOT_11
timestamp 1355475633
transform 0 1 951 -1 0 -234
box -5 -23 43 41
use NOT  NOT_3
timestamp 1355475633
transform 0 1 1152 -1 0 -212
box -5 -23 43 41
use NOT  NOT_4
timestamp 1355475633
transform 0 1 1152 -1 0 -240
box -5 -23 43 41
use NOR  NOR_1
timestamp 1355475848
transform 0 1 262 -1 0 -304
box -14 -22 34 42
use NOT  NOT_10
timestamp 1355475633
transform 0 1 785 -1 0 -290
box -5 -23 43 41
use NOT  NOT_5
timestamp 1355475633
transform 0 1 1152 -1 0 -268
box -5 -23 43 41
use NOT  NOT_7
timestamp 1355475633
transform 0 1 263 -1 0 -343
box -5 -23 43 41
use NAND  NAND_6
timestamp 1355475793
transform 0 1 767 -1 0 -355
box -16 -2 32 62
<< labels >>
rlabel space 28 63 28 63 5 Vdd
rlabel space 12 41 12 41 3 In1
rlabel space 12 33 12 33 3 In2
rlabel m2contact 12 27 12 27 3 S
rlabel metal2 158 38 158 38 1 Clkb
rlabel metal2 169 31 169 31 1 Clk
rlabel space 413 21 417 22 1 ClkB
rlabel space 713 21 717 22 1 ClkB
rlabel space 822 21 826 22 1 ClkB
rlabel space 835 21 839 22 1 RstB
rlabel m2contact 918 -53 922 -49 1 GO?
rlabel space 1059 21 1063 22 1 ClkB
rlabel metal1 1160 -292 1160 -292 5 In
rlabel metal1 1187 -300 1187 -300 3 pos
rlabel metal1 1135 -299 1135 -299 3 Vneg
rlabel space 15 5 15 5 1 Gnd
rlabel m2contact 1160 -395 1160 -395 1 Out
rlabel metal2 150 -429 151 -428 1 RST_IR
rlabel metal2 271 -425 271 -425 1 DIS_CO?
rlabel metal2 392 -428 392 -428 1 Iin?
rlabel metal2 469 -428 469 -427 1 MSB_CE
rlabel metal2 544 -428 544 -428 1 C1?
rlabel metal2 622 -426 622 -426 1 C2?
rlabel metal2 728 -427 728 -427 1 RST_C2_C0?
rlabel metal2 797 -428 797 -428 1 RST_C1_CO?
rlabel metal2 875 -426 875 -426 1 LSB_CE
rlabel metal2 960 -426 960 -425 1 C2Ref?
rlabel metal2 1160 -429 1160 -429 1 W_OUT
<< end >>
