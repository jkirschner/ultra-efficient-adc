* SPICE3 file created from msb_registers.ext - technology: scmos

.subckt ToggleFlipFlop_Low_Layout ClkB Vpos Qb Vneg RstB Q Clk T
M1000 a_177_n338# T Vpos Vpos pfet w=6u l=0.9u
+ ad=9p pd=15u as=189.36p ps=301.8u 
M1001 a_194_n255# a_177_n289# Vpos Vpos pfet w=6u l=0.9u
+ ad=18p pd=18u as=0p ps=0u 
M1002 Vpos a_195_n289# a_194_n255# Vpos pfet w=6u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1003 a_227_n262# RstB Vpos Vpos pfet w=12.6u l=0.9u
+ ad=44.28p pd=64.2u as=0p ps=0u 
M1004 Vpos RstB a_227_n262# Vpos pfet w=7.8u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1005 a_227_n262# RstB Vpos Vpos pfet w=7.8u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1006 Vpos RstB a_227_n262# Vpos pfet w=7.8u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1007 Vpos a_227_n262# a_225_n326# Vpos pfet w=6u l=0.9u
+ ad=0p pd=0u as=6.66p ps=15u 
M1008 a_266_n262# RstB Vpos Vpos pfet w=12.6u l=0.9u
+ ad=44.28p pd=64.2u as=0p ps=0u 
M1009 Vpos RstB a_266_n262# Vpos pfet w=7.8u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1010 a_266_n262# RstB Vpos Vpos pfet w=7.8u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1011 Vpos RstB a_266_n262# Vpos pfet w=7.8u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1012 Vpos a_266_n262# a_258_n330# Vpos pfet w=6u l=0.9u
+ ad=0p pd=0u as=6.12p ps=15u 
M1013 a_177_n289# T Vpos Vpos pfet w=6u l=0.9u
+ ad=10.8p pd=15.6u as=0p ps=0u 
M1014 Vpos Q a_177_n289# Vpos pfet w=6u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1015 a_195_n289# a_177_n338# Vpos Vpos pfet w=6u l=0.9u
+ ad=10.8p pd=15.6u as=0p ps=0u 
M1016 Vpos Qb a_195_n289# Vpos pfet w=6u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1017 a_229_n289# a_194_n255# Vpos Vpos pfet w=6u l=0.9u
+ ad=7.2p pd=14.4u as=0p ps=0u 
M1018 a_227_n262# ClkB a_229_n289# Vpos pfet w=6u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1019 a_245_n289# Clk a_227_n262# Vpos pfet w=6u l=0.9u
+ ad=7.2p pd=14.4u as=0p ps=0u 
M1020 Vpos a_225_n326# a_245_n289# Vpos pfet w=6u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1021 a_261_n289# a_225_n326# Vpos Vpos pfet w=6u l=0.9u
+ ad=7.2p pd=14.4u as=0p ps=0u 
M1022 a_266_n262# Clk a_261_n289# Vpos pfet w=6u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1023 a_277_n289# ClkB a_266_n262# Vpos pfet w=6u l=0.9u
+ ad=7.2p pd=14.4u as=0p ps=0u 
M1024 Vpos a_258_n330# a_277_n289# Vpos pfet w=6u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1025 a_172_n313# T Vneg Vneg nfet w=3u l=0.9u
+ ad=5.4p pd=9.6u as=48.96p ps=94.8u 
M1026 a_177_n289# Q a_172_n313# Vneg nfet w=3u l=0.9u
+ ad=4.5p pd=9u as=0p ps=0u 
M1027 a_198_n313# a_177_n338# Vneg Vneg nfet w=3u l=0.9u
+ ad=2.7p pd=7.8u as=0p ps=0u 
M1028 a_195_n289# Qb a_198_n313# Vneg nfet w=3u l=0.9u
+ ad=4.5p pd=9u as=0p ps=0u 
M1029 Qb a_258_n330# Vpos Vpos pfet w=6u l=0.9u
+ ad=7.29p pd=15.6u as=0p ps=0u 
M1030 Q a_266_n262# Vpos Vpos pfet w=6u l=0.9u
+ ad=8.64p pd=15u as=0p ps=0u 
M1031 a_229_n320# a_225_n326# Vneg Vneg nfet w=3u l=0.9u
+ ad=3.6p pd=8.4u as=0p ps=0u 
M1032 a_227_n262# ClkB a_229_n320# Vneg nfet w=3u l=0.9u
+ ad=5.4p pd=9.6u as=0p ps=0u 
M1033 a_245_n320# Clk a_227_n262# Vneg nfet w=3u l=0.9u
+ ad=3.6p pd=8.4u as=0p ps=0u 
M1034 Vneg a_194_n255# a_245_n320# Vneg nfet w=3u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1035 a_261_n320# a_258_n330# Vneg Vneg nfet w=3u l=0.9u
+ ad=3.6p pd=8.4u as=0p ps=0u 
M1036 a_266_n262# Clk a_261_n320# Vneg nfet w=3u l=0.9u
+ ad=5.4p pd=9.6u as=0p ps=0u 
M1037 a_277_n320# ClkB a_266_n262# Vneg nfet w=3u l=0.9u
+ ad=3.6p pd=8.4u as=0p ps=0u 
M1038 Vneg a_225_n326# a_277_n320# Vneg nfet w=3u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1039 Qb a_258_n330# Vneg Vneg nfet w=3u l=0.9u
+ ad=5.4p pd=9.6u as=0p ps=0u 
M1040 a_177_n338# T Vneg Vneg nfet w=3u l=0.9u
+ ad=5.4p pd=9.6u as=0p ps=0u 
M1041 a_195_n338# a_177_n289# Vneg Vneg nfet w=3u l=0.9u
+ ad=5.4p pd=9.6u as=0p ps=0u 
M1042 a_194_n255# a_195_n289# a_195_n338# Vneg nfet w=3u l=0.9u
+ ad=3.78p pd=9u as=0p ps=0u 
M1043 a_225_n326# a_227_n262# Vneg Vneg nfet w=3u l=0.9u
+ ad=4.5p pd=9u as=0p ps=0u 
M1044 a_258_n330# a_266_n262# Vneg Vneg nfet w=3u l=0.9u
+ ad=4.5p pd=9u as=0p ps=0u 
M1045 Q a_266_n262# Vneg Vneg nfet w=3u l=0.9u
+ ad=4.23p pd=9u as=0p ps=0u 
.ends

.subckt ResetFlipFlop_Low_Layout ClkB Vpos D Vneg RstB Q Clk
M1000 a_227_n262# RstB Vpos Vpos pfet w=12.6u l=0.9u
+ ad=44.28p pd=64.2u as=135.54p ps=211.2u 
M1001 Vpos RstB a_227_n262# Vpos pfet w=7.8u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1002 a_227_n262# RstB Vpos Vpos pfet w=7.8u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1003 Vpos RstB a_227_n262# Vpos pfet w=7.8u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1004 Vpos a_227_n262# a_225_n326# Vpos pfet w=6u l=0.9u
+ ad=0p pd=0u as=6.66p ps=15u 
M1005 a_266_n262# RstB Vpos Vpos pfet w=12.6u l=0.9u
+ ad=44.28p pd=64.2u as=0p ps=0u 
M1006 Vpos RstB a_266_n262# Vpos pfet w=7.8u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1007 a_266_n262# RstB Vpos Vpos pfet w=7.8u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1008 Vpos RstB a_266_n262# Vpos pfet w=7.8u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1009 Vpos a_266_n262# a_258_n330# Vpos pfet w=6u l=0.9u
+ ad=0p pd=0u as=6.12p ps=15u 
M1010 a_229_n289# D Vpos Vpos pfet w=6u l=0.9u
+ ad=7.2p pd=14.4u as=0p ps=0u 
M1011 a_227_n262# ClkB a_229_n289# Vpos pfet w=6u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1012 a_245_n289# Clk a_227_n262# Vpos pfet w=6u l=0.9u
+ ad=7.2p pd=14.4u as=0p ps=0u 
M1013 Vpos a_225_n326# a_245_n289# Vpos pfet w=6u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1014 a_261_n289# a_225_n326# Vpos Vpos pfet w=6u l=0.9u
+ ad=7.2p pd=14.4u as=0p ps=0u 
M1015 a_266_n262# Clk a_261_n289# Vpos pfet w=6u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1016 a_277_n289# ClkB a_266_n262# Vpos pfet w=6u l=0.9u
+ ad=7.2p pd=14.4u as=0p ps=0u 
M1017 Vpos a_258_n330# a_277_n289# Vpos pfet w=6u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1018 Qb a_258_n330# Vpos Vpos pfet w=6u l=0.9u
+ ad=7.29p pd=15.6u as=0p ps=0u 
M1019 Q a_266_n262# Vpos Vpos pfet w=6u l=0.9u
+ ad=8.64p pd=15u as=0p ps=0u 
M1020 a_229_n320# a_225_n326# Vneg Vneg nfet w=3u l=0.9u
+ ad=3.6p pd=8.4u as=30.96p ps=58.8u 
M1021 a_227_n262# ClkB a_229_n320# Vneg nfet w=3u l=0.9u
+ ad=5.4p pd=9.6u as=0p ps=0u 
M1022 a_245_n320# Clk a_227_n262# Vneg nfet w=3u l=0.9u
+ ad=3.6p pd=8.4u as=0p ps=0u 
M1023 Vneg D a_245_n320# Vneg nfet w=3u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1024 a_261_n320# a_258_n330# Vneg Vneg nfet w=3u l=0.9u
+ ad=3.6p pd=8.4u as=0p ps=0u 
M1025 a_266_n262# Clk a_261_n320# Vneg nfet w=3u l=0.9u
+ ad=5.4p pd=9.6u as=0p ps=0u 
M1026 a_277_n320# ClkB a_266_n262# Vneg nfet w=3u l=0.9u
+ ad=3.6p pd=8.4u as=0p ps=0u 
M1027 Vneg a_225_n326# a_277_n320# Vneg nfet w=3u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1028 Qb a_258_n330# Vneg Vneg nfet w=3u l=0.9u
+ ad=5.4p pd=9.6u as=0p ps=0u 
M1029 a_225_n326# a_227_n262# Vneg Vneg nfet w=3u l=0.9u
+ ad=4.5p pd=9u as=0p ps=0u 
M1030 a_258_n330# a_266_n262# Vneg Vneg nfet w=3u l=0.9u
+ ad=4.5p pd=9u as=0p ps=0u 
M1031 Q a_266_n262# Vneg Vneg nfet w=3u l=0.9u
+ ad=4.23p pd=9u as=0p ps=0u 
.ends


* Top level circuit msb_registers

X0 ToggleFlipFlop_Low_Layout_1/Qb pos ToggleFlipFlop_Low_Layout_0/Qb neg RST_IRb ResetFlipFlop_Low_Layout_1/D ResetFlipFlop_Low_Layout_0/D MSB_CLK ToggleFlipFlop_Low_Layout
X1 SYS_CLKb pos ToggleFlipFlop_Low_Layout_1/Qb neg RST_IRb ResetFlipFlop_Low_Layout_0/D SYS_CLK MSB_CLK ToggleFlipFlop_Low_Layout
X2 W_CLKb pos ResetFlipFlop_Low_Layout_1/D neg RST_ORb Bit0 W_CLK ResetFlipFlop_Low_Layout
X3 W_CLKb pos ResetFlipFlop_Low_Layout_0/D neg RST_ORb Bit1 W_CLK ResetFlipFlop_Low_Layout
.end

