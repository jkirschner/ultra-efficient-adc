magic
tech scmos
timestamp 1355475992
<< nwell >>
rect -12 -11 36 26
<< pwell >>
rect -12 -42 36 -11
<< ntransistor >>
rect 0 -31 3 -21
rect 9 -31 12 -21
rect 18 -31 21 -21
<< ptransistor >>
rect 0 0 3 20
rect 9 0 12 20
rect 18 0 21 20
<< ndiffusion >>
rect -3 -27 0 -21
rect -1 -31 0 -27
rect 3 -31 9 -21
rect 12 -31 18 -21
rect 21 -22 24 -21
rect 21 -26 22 -22
rect 21 -31 24 -26
<< pdiffusion >>
rect -3 19 0 20
rect -1 15 0 19
rect -3 0 0 15
rect 3 6 9 20
rect 3 2 4 6
rect 8 2 9 6
rect 3 0 9 2
rect 12 19 18 20
rect 12 15 13 19
rect 17 15 18 19
rect 12 0 18 15
rect 21 6 24 20
rect 21 2 22 6
rect 21 0 24 2
<< ndcontact >>
rect -5 -31 -1 -27
rect 22 -26 26 -22
<< pdcontact >>
rect -5 15 -1 19
rect 4 2 8 6
rect 13 15 17 19
rect 22 2 26 6
<< psubstratepcontact >>
rect 21 -39 25 -35
<< nsubstratencontact >>
rect 28 15 32 19
<< polysilicon >>
rect 0 20 3 22
rect 9 20 12 22
rect 18 20 21 22
rect 0 -1 3 0
rect 0 -21 3 -5
rect 9 -8 12 0
rect 9 -21 12 -12
rect 18 -15 21 0
rect 18 -21 21 -19
rect 0 -33 3 -31
rect 9 -33 12 -31
rect 18 -33 21 -31
<< polycontact >>
rect -1 -5 3 -1
rect 8 -12 12 -8
rect 17 -19 21 -15
<< metal1 >>
rect -11 19 36 22
rect -11 15 -5 19
rect -1 15 13 19
rect 17 15 28 19
rect 32 15 36 19
rect -11 9 36 15
rect 8 2 22 6
rect 26 2 28 6
rect -12 -5 -1 -1
rect 24 -8 28 2
rect -12 -12 8 -8
rect 24 -12 36 -8
rect -12 -19 17 -15
rect 24 -22 28 -12
rect 26 -26 28 -22
rect -12 -31 -5 -29
rect -1 -31 36 -29
rect -12 -35 36 -31
rect -12 -39 21 -35
rect 25 -39 36 -35
rect -12 -42 36 -39
<< labels >>
rlabel metal1 34 -10 35 -10 7 Out
rlabel metal1 -11 -3 -11 -3 3 A
rlabel metal1 -11 -10 -11 -10 3 B
rlabel metal1 -11 -17 -11 -17 3 C
rlabel metal1 -3 -39 -3 -39 1 neg
rlabel metal1 -8 16 -8 16 3 pos
<< end >>
