magic
tech scmos
timestamp 1355723001
<< nwell >>
rect -1243 3082 -1239 3103
<< pwell >>
rect -868 2952 -864 2963
rect -1067 2931 -997 2936
rect -273 2903 -265 2914
rect -273 2897 -235 2903
<< electrodecap >>
rect -1232 2096 -1227 2101
<< polysilicon >>
rect -1232 2096 -1227 2101
<< metal1 >>
rect -1273 3107 -1251 3216
rect -977 3111 -905 3121
rect -1243 3082 -1239 3099
rect -1029 3097 -1019 3101
rect -978 3097 -949 3101
rect -1029 3076 -1025 3097
rect -914 3076 -905 3111
rect -218 3113 -204 3216
rect -218 3109 -214 3113
rect -206 3109 -204 3113
rect -193 3195 -176 3217
rect -193 3184 379 3195
rect -193 3095 -183 3184
rect -914 3072 -909 3076
rect 128 3039 144 3056
rect 128 3001 151 3039
rect -135 2903 -100 2918
rect -265 2902 -235 2903
rect -265 2899 -222 2902
rect -273 2897 -222 2899
rect -1303 2775 -1141 2795
rect -1303 2774 -1205 2775
rect -1149 2774 -1141 2775
rect -1303 2650 -1281 2774
rect -248 2683 -222 2897
rect 196 2740 209 3123
rect 369 3107 379 3184
rect 357 3086 379 3107
rect 196 2726 197 2740
rect 226 2690 242 2894
rect 164 2661 200 2665
rect -1303 2444 -1280 2650
rect -1303 2431 -1288 2444
rect -1282 2431 -1280 2444
rect -1303 2204 -1280 2431
rect -1261 2628 -1169 2652
rect -1140 2647 -1122 2654
rect -1261 2501 -1226 2628
rect -787 2604 3 2619
rect 169 2592 222 2597
rect -1261 2490 -1149 2501
rect -1261 2231 -1226 2490
rect -1167 2479 -1149 2490
rect -310 2442 -300 2574
rect -248 2454 -222 2574
rect -101 2571 328 2575
rect 336 2514 360 2582
rect 377 2575 381 2582
rect 374 2571 381 2575
rect 377 2522 381 2571
rect 386 2531 391 2581
rect 386 2525 463 2531
rect 377 2517 436 2522
rect 336 2494 410 2514
rect -248 2429 -66 2454
rect -997 2396 -409 2397
rect -1184 2375 -1180 2395
rect -992 2384 -409 2396
rect -992 2383 -393 2384
rect -992 2382 -981 2383
rect -1184 2363 -212 2375
rect -1191 2352 -473 2353
rect -1180 2342 -473 2352
rect -1180 2341 -462 2342
rect -1180 2314 -542 2325
rect -1108 2301 -11 2302
rect -1108 2289 10 2301
rect -1118 2288 10 2289
rect -968 2276 -724 2282
rect -461 2266 -27 2279
rect -782 2248 -590 2257
rect -1303 2179 -1258 2204
rect -600 2189 -590 2248
rect -461 2245 -450 2266
rect -494 2237 -450 2245
rect -582 2217 -559 2221
rect -555 2202 -551 2207
rect -600 2177 -557 2189
rect -782 2152 -564 2156
rect -782 2142 -778 2152
rect -582 2145 -559 2149
rect -461 2129 -450 2237
rect -319 2214 -300 2266
rect -173 2192 -90 2201
rect -494 2121 -450 2129
rect -379 2145 -373 2152
rect -364 2145 -363 2152
rect -1316 1728 -390 1745
rect -1316 1706 -390 1723
rect -379 -80 -363 2145
rect -182 2059 -142 2074
rect -103 1833 -90 2192
rect -141 1816 -90 1833
rect -66 2093 -50 2097
rect -308 1784 -304 1797
rect -289 1424 -238 1445
rect -289 -86 -255 1424
rect -141 1339 -124 1816
rect -66 1577 -50 2081
rect -8 1597 10 2288
rect 177 1953 185 2133
rect 300 1611 301 1622
rect 305 1611 306 1622
rect -88 1565 -50 1577
rect -88 1447 -72 1565
rect 259 1563 274 1611
rect 300 1607 306 1611
rect 300 1563 306 1566
rect 325 1564 348 1611
rect 300 1552 301 1563
rect 305 1552 306 1563
rect 392 1529 400 1684
rect 418 1622 436 2517
rect 423 1611 436 1622
rect 418 1563 436 1611
rect 406 1554 436 1563
rect 406 1529 414 1554
rect -12 1507 4 1512
rect 445 1511 463 2525
rect -88 1432 -33 1447
rect -140 -85 -124 1339
rect -53 -61 -33 1432
rect 19 -9 37 19
rect 48 0 79 7
rect 48 -8 52 0
rect 129 -7 152 16
rect 65 -17 152 -7
rect 47 -52 49 -51
rect 50 -52 52 -51
rect 47 -61 52 -52
rect -53 -76 52 -61
rect 235 -76 262 76
<< m2contact >>
rect -1243 3099 -1239 3103
rect -1029 3072 -1025 3076
rect -214 3109 -206 3113
rect 196 3123 209 3142
rect -909 3072 -905 3076
rect -81 3039 -74 3056
rect 144 3039 151 3056
rect -880 3014 -872 3018
rect -771 3003 -767 3018
rect -581 3004 -573 3008
rect -470 3004 -462 3008
rect -362 3004 -354 3008
rect -868 2952 -864 2963
rect -273 2899 -265 2904
rect -100 2903 -95 2918
rect 14 2904 18 2918
rect 197 2726 209 2740
rect -248 2671 -222 2683
rect 159 2661 164 2665
rect 238 2661 243 2665
rect -1288 2431 -1282 2444
rect -798 2604 -787 2619
rect 3 2603 9 2619
rect 222 2590 230 2597
rect -310 2574 -300 2583
rect -1186 2472 -1180 2482
rect -1211 2431 -1205 2444
rect -1185 2433 -1178 2441
rect -310 2429 -300 2442
rect -248 2574 -222 2583
rect 18 2580 45 2587
rect -107 2571 -101 2575
rect 328 2571 332 2575
rect 368 2580 373 2584
rect 370 2571 374 2575
rect 19 2504 46 2511
rect 70 2482 87 2494
rect -66 2429 -49 2454
rect -1001 2382 -992 2396
rect -409 2384 -393 2397
rect -212 2363 -197 2375
rect -1191 2341 -1180 2352
rect -473 2342 -462 2353
rect -1190 2314 -1180 2325
rect -542 2314 -530 2325
rect -1118 2289 -1108 2302
rect -974 2276 -968 2282
rect -724 2275 -717 2283
rect -1271 2214 -1263 2219
rect -587 2217 -582 2221
rect -563 2210 -559 2214
rect -564 2152 -559 2156
rect -587 2145 -582 2149
rect -783 2126 -779 2130
rect -27 2265 -16 2279
rect -373 2145 -364 2152
rect -390 1728 -385 1745
rect -390 1706 -385 1723
rect -142 2059 -130 2074
rect -207 1822 -201 1830
rect -66 2081 -50 2093
rect -308 1780 -304 1784
rect 19 2265 28 2279
rect 177 2133 185 2140
rect 129 2060 151 2074
rect 382 1684 400 1701
rect 301 1611 305 1622
rect 301 1552 305 1563
rect -13 1521 -8 1540
rect 19 1521 24 1540
rect 418 1611 423 1622
rect -56 1507 -51 1512
rect 177 1501 185 1511
rect 445 1499 463 1511
rect -12 1487 -8 1494
rect 146 1487 152 1494
<< metal2 >>
rect -451 3142 -426 3216
rect 437 3149 518 3165
rect -1243 3123 196 3142
rect -1243 3103 -1236 3123
rect -1239 3099 -1236 3103
rect -1300 3089 -1246 3094
rect -1300 2843 -1287 3089
rect -1025 3072 -987 3076
rect -992 3006 -987 3072
rect -909 3069 -905 3072
rect -909 3065 -864 3069
rect -1001 3001 -987 3006
rect -1001 2936 -997 3001
rect -868 2963 -864 3065
rect -74 3039 144 3056
rect 437 3008 518 3024
rect -280 3003 -266 3007
rect -1067 2931 -997 2936
rect -273 2914 -266 3003
rect -273 2904 -265 2914
rect -95 2904 14 2918
rect -95 2903 8 2904
rect -1300 2835 -1178 2843
rect -1189 2482 -1178 2835
rect 180 2740 209 2741
rect 180 2726 197 2740
rect -1189 2472 -1186 2482
rect -1180 2472 -1178 2482
rect -1282 2431 -1211 2444
rect -1178 2433 -1133 2441
rect -1291 2341 -1191 2352
rect -1180 2341 -1179 2352
rect -1291 2151 -1280 2341
rect -1271 2314 -1190 2325
rect -1271 2219 -1263 2314
rect -1142 2295 -1133 2433
rect -1183 2287 -1133 2295
rect -1118 2302 -1108 2624
rect -1000 2413 -991 2627
rect -1000 2396 -992 2413
rect -1183 2253 -1178 2287
rect -1118 2244 -1108 2289
rect -974 2282 -968 2283
rect -997 2256 -993 2267
rect -974 2257 -968 2276
rect -881 2271 -872 2622
rect -725 2283 -717 2626
rect -725 2275 -724 2283
rect -965 2262 -872 2271
rect -646 2267 -638 2626
rect -542 2325 -530 2626
rect -473 2353 -462 2627
rect -392 2495 -386 2625
rect -310 2583 -300 2627
rect -248 2583 -222 2671
rect 179 2661 238 2665
rect -107 2575 -101 2625
rect 3 2619 9 2628
rect 18 2511 45 2580
rect 18 2504 19 2511
rect 158 2509 164 2581
rect 179 2514 184 2582
rect 171 2509 184 2514
rect -392 2494 87 2495
rect -392 2482 70 2494
rect -436 2441 -310 2442
rect -437 2429 -310 2441
rect -437 2281 -427 2429
rect -965 2254 -957 2262
rect -837 2259 -638 2267
rect -587 2274 -427 2281
rect -393 2384 -392 2397
rect -837 2241 -829 2259
rect -837 2233 -828 2241
rect -587 2221 -582 2274
rect -409 2242 -392 2384
rect -212 2250 -197 2363
rect -409 2234 -331 2242
rect -335 2229 -331 2234
rect -1291 2140 -1266 2151
rect -587 2149 -582 2217
rect -579 2210 -563 2214
rect -579 2136 -574 2210
rect -506 2208 -395 2217
rect -571 2202 -550 2207
rect -571 2156 -566 2202
rect -571 2152 -564 2156
rect -496 2144 -425 2153
rect -555 2136 -551 2144
rect -579 2131 -551 2136
rect -579 2130 -574 2131
rect -779 2126 -574 2130
rect -433 1688 -425 2144
rect -403 1700 -395 2208
rect -364 2147 -360 2151
rect -66 2093 -50 2429
rect -16 2265 19 2279
rect 222 2140 230 2590
rect 373 2580 385 2584
rect 332 2571 370 2575
rect 381 2517 385 2580
rect 185 2133 230 2140
rect -130 2060 129 2074
rect 151 2060 152 2074
rect -351 1780 -308 1784
rect -351 1774 -304 1780
rect -351 1745 -343 1774
rect -385 1728 -343 1745
rect -298 1723 -294 1732
rect -385 1706 -294 1723
rect 368 1701 385 2517
rect -403 1692 -342 1700
rect -396 1691 -342 1692
rect -433 1679 -342 1688
rect 368 1684 382 1701
rect -433 1677 -425 1679
rect 305 1611 418 1622
rect 305 1552 386 1563
rect -8 1521 19 1540
rect 378 1512 386 1552
rect -51 1511 185 1512
rect -51 1507 177 1511
rect -56 1502 177 1507
rect 378 1511 463 1512
rect 378 1499 445 1511
rect -8 1487 146 1494
rect 416 1399 497 1415
rect 419 1249 500 1265
rect 419 1101 500 1117
rect 418 952 499 968
rect 418 802 499 818
rect 419 651 500 667
rect 418 501 499 517
rect 418 352 499 368
rect 417 203 498 219
rect 418 53 499 69
<< pseudo_rmetal2 >>
rect -872 3018 -870 3022
<< m3contact >>
rect -1003 3020 -999 3024
rect -880 3018 -872 3022
rect -767 3003 -763 3018
rect -581 3008 -573 3012
rect -470 3008 -462 3012
rect -362 3008 -354 3012
rect -997 2267 -992 2272
rect -1005 2256 -1000 2261
rect -201 1822 -195 1830
<< metal3 >>
rect -1033 3065 -1023 3216
rect -1033 3057 -996 3065
rect -1004 3024 -996 3057
rect -1004 3020 -1003 3024
rect -999 3020 -996 3024
rect -1004 3019 -996 3020
rect -881 3022 -871 3216
rect -881 3018 -880 3022
rect -872 3018 -871 3022
rect -881 3017 -871 3018
rect -772 3018 -762 3216
rect -772 3012 -767 3018
rect -768 3003 -767 3012
rect -763 3003 -762 3018
rect -582 3012 -572 3216
rect -582 3008 -581 3012
rect -573 3008 -572 3012
rect -582 3007 -572 3008
rect -471 3012 -461 3216
rect -362 3021 -353 3216
rect -471 3008 -470 3012
rect -462 3008 -461 3012
rect -471 3007 -461 3008
rect -363 3012 -353 3021
rect -363 3008 -362 3012
rect -354 3008 -353 3012
rect -363 3007 -353 3008
rect -768 3002 -762 3003
rect 398 2551 416 3217
rect -128 2534 416 2551
rect -1328 2272 -991 2279
rect -1328 2268 -997 2272
rect -998 2267 -997 2268
rect -992 2267 -991 2272
rect -998 2266 -991 2267
rect -1328 2261 -999 2262
rect -1328 2256 -1005 2261
rect -1000 2256 -999 2261
rect -1328 2251 -999 2256
rect -128 1896 -114 2534
rect -155 1884 -114 1896
rect -155 1831 -144 1884
rect -202 1830 -144 1831
rect -202 1822 -201 1830
rect -195 1822 -144 1830
rect -202 1821 -144 1822
use NOT  NOT_4
timestamp 1355475633
transform -1 0 -978 0 -1 3107
box -5 -23 43 41
use stateMachine  stateMachine_0
timestamp 1355540337
transform 1 0 -1265 0 1 3050
box -14 -441 1196 68
use NOT  NOT_3
timestamp 1355475633
transform -1 0 238 0 -1 2671
box -5 -23 43 41
use msb_registers  msb_registers_0
timestamp 1355455137
transform 0 1 227 1 0 2875
box -295 -224 301 222
use NOT  NOT_6
timestamp 1355475633
transform 0 1 -1190 1 0 2439
box -5 -23 43 41
use NOT  NOT_5
timestamp 1355475633
transform 0 1 -1190 1 0 2395
box -5 -23 43 41
use SPDT  SPDT_0
timestamp 1355531441
transform 1 0 -597 0 -1 2246
box 38 1 105 68
use SPDT  SPDT_1
timestamp 1355531441
transform 1 0 -597 0 1 2120
box 38 1 105 68
use AnalogSwitch  AnalogSwitch_0
timestamp 1355620377
transform 1 0 -944 0 1 2213
box -325 -461 424 47
use Comparator  Comparator_0
timestamp 1355695794
transform 0 1 -336 1 0 1439
box -6 -28 815 195
use NOT  NOT_2
timestamp 1355475633
transform 0 1 295 -1 0 1606
box -5 -23 43 41
use NOT  NOT_1
timestamp 1355475633
transform -1 0 -13 0 -1 1517
box -5 -23 43 41
use lsb_registers_Layout  lsb_registers_Layout_0
timestamp 1355674588
transform 0 1 263 -1 0 1521
box -990 -263 1521 160
use NOT  NOT_0
timestamp 1355475633
transform 0 1 42 -1 0 -12
box -5 -23 43 41
<< labels >>
rlabel metal1 49 -72 49 -72 1 GO?
rlabel metal2 -1240 3124 -1240 3124 1 CLK
rlabel metal2 490 1405 490 1405 1 Bit11
rlabel metal2 492 60 492 60 1 Bit2
rlabel metal2 492 211 492 211 1 Bit3
rlabel metal2 493 359 493 359 1 Bit4
rlabel metal2 488 508 488 508 1 Bit5
rlabel metal2 490 659 490 659 1 Bit6
rlabel metal2 491 809 491 809 1 Bit7
rlabel metal2 486 959 486 959 1 Bit8
rlabel metal2 488 1108 488 1108 1 Bit9
rlabel metal2 490 1256 490 1256 1 Bit10
rlabel metal2 500 3157 500 3157 1 Bit0
rlabel metal2 503 3014 503 3014 1 Bit1
rlabel metal1 -371 -74 -371 -74 1 Vpw1
rlabel metal1 -133 -77 -133 -77 1 Vpw2
rlabel metal1 -273 -76 -273 -76 1 Bias
rlabel metal2 -437 3208 -437 3208 1 CLK
rlabel metal2 -433 2151 -433 2151 1 Comp_Vthresh
rlabel metal2 -433 2215 -433 2215 1 Comp_Vin
rlabel metal1 -1308 1714 -1308 1714 1 V-
rlabel metal1 -1308 1737 -1308 1737 1 V+
rlabel metal1 -211 3211 -211 3211 1 Sexit
rlabel metal3 -358 3210 -358 3210 1 S2x
rlabel metal3 -466 3211 -466 3211 1 Svt
rlabel metal3 -578 3211 -578 3211 1 Stv
rlabel metal3 -767 3212 -767 3212 1 Sref
rlabel metal3 -876 3211 -876 3211 1 Sin
rlabel metal3 -1028 3210 -1028 3210 1 Sreset
rlabel metal3 -1319 2272 -1319 2272 1 Iin
rlabel metal3 -1319 2256 -1319 2256 1 Iref
rlabel metal1 -185 3212 -185 3212 5 RSTb
rlabel metal3 409 3205 409 3205 1 PosA
rlabel metal1 249 -68 249 -68 1 Vneg
rlabel metal1 -1261 3207 -1261 3207 1 Vpos
<< end >>
