* SPICE3 file created from GainLatch_layout.ext - technology: scmos

M1000 a_26_61# Cascode N1 PosA pfet w=4.8u l=2.4u
+ ad=29.52p pd=43.2u as=27p ps=46.8u 
M1001 PosA Vbias a_26_61# PosA pfet w=9u l=18u
+ ad=16.2p pd=21.6u as=0p ps=0u 
M1002 a_26_61# Vbias PosA PosA pfet w=9u l=18u
+ ad=0p pd=0u as=0p ps=0u 
M1003 N1 Cascode a_26_61# PosA pfet w=4.8u l=2.4u
+ ad=0p pd=0u as=0p ps=0u 
M1004 PosD a_22_4# a_19_27# PosA pfet w=4.5u l=2.7u
+ ad=16.2p pd=25.2u as=15.48p ps=34.8u 
M1005 a_33_11# a_33_11# PosD PosA pfet w=4.5u l=2.7u
+ ad=13.5p pd=24u as=0p ps=0u 
M1006 N1 Vp N3 PosA pfet w=3.6u l=3.6u
+ ad=0p pd=0u as=10.8p ps=20.4u 
M1007 N2 a_80_23# N1 PosA pfet w=3.6u l=3.6u
+ ad=6.48p pd=10.8u as=0p ps=0u 
M1008 N1 a_80_23# N2 PosA pfet w=3.6u l=3.6u
+ ad=0p pd=0u as=0p ps=0u 
M1009 N3 Vp N1 PosA pfet w=3.6u l=3.6u
+ ad=0p pd=0u as=0p ps=0u 
M1010 PosD a_33_11# a_33_11# PosA pfet w=4.5u l=2.7u
+ ad=0p pd=0u as=0p ps=0u 
M1011 a_19_27# a_22_4# PosD PosA pfet w=4.5u l=2.7u
+ ad=0p pd=0u as=0p ps=0u 
M1012 a_35_n9# a_33_11# a_19_27# PosA pfet w=0.9u l=0.6u
+ ad=3.42p pd=10.8u as=0p ps=0u 
M1013 a_19_27# a_33_11# a_35_n9# PosA pfet w=0.9u l=0.6u
+ ad=0p pd=0u as=0p ps=0u 
M1014 a_35_n9# a_22_4# Vneg Vneg nfet w=3.6u l=1.8u
+ ad=16.92p pd=36u as=36.72p ps=74.4u 
M1015 Vneg N3 a_35_n9# Vneg nfet w=2.4u l=2.7u
+ ad=0p pd=0u as=0p ps=0u 
M1016 N3 N3 Vneg Vneg nfet w=2.4u l=2.7u
+ ad=4.32p pd=8.4u as=0p ps=0u 
M1017 Vneg N3 N3 Vneg nfet w=2.4u l=2.7u
+ ad=0p pd=0u as=0p ps=0u 
M1018 a_35_n9# N3 Vneg Vneg nfet w=2.4u l=2.7u
+ ad=0p pd=0u as=0p ps=0u 
M1019 Vneg a_22_4# a_35_n9# Vneg nfet w=3.6u l=1.8u
+ ad=0p pd=0u as=0p ps=0u 
M1020 a_33_11# a_35_n9# Vneg Vneg nfet w=3.6u l=1.8u
+ ad=16.92p pd=36u as=0p ps=0u 
M1021 Vneg N2 a_33_11# Vneg nfet w=2.4u l=2.7u
+ ad=0p pd=0u as=0p ps=0u 
M1022 N2 N2 Vneg Vneg nfet w=2.4u l=2.7u
+ ad=4.32p pd=8.4u as=0p ps=0u 
M1023 Vneg N2 N2 Vneg nfet w=2.4u l=2.7u
+ ad=0p pd=0u as=0p ps=0u 
M1024 a_33_11# N2 Vneg Vneg nfet w=2.4u l=2.7u
+ ad=0p pd=0u as=0p ps=0u 
M1025 Vneg a_35_n9# a_33_11# Vneg nfet w=3.6u l=1.8u
+ ad=0p pd=0u as=0p ps=0u 
