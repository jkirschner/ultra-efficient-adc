magic
tech scmos
timestamp 1355692754
<< end >>
