magic
tech scmos
timestamp 1355184513
<< electrodecontact >>
rect 11 -117 15 -113
rect 86 -115 90 -111
<< electrodecap >>
rect -292 -456 57 -107
rect 70 -456 419 -107
<< ntransistor >>
rect -8 -23 -5 -13
rect 1 -23 4 -13
rect 10 -23 13 -13
rect 19 -23 22 -13
rect 36 -23 39 -13
rect 43 -23 46 -13
rect 61 -23 64 -13
rect 78 -23 81 -13
rect 87 -23 90 -13
rect 104 -23 107 -13
rect 113 -23 116 -13
rect 130 -23 133 -13
rect 139 -23 142 -13
rect 8 -95 10 -71
rect 83 -89 85 -65
<< ptransistor >>
rect -8 -1 -5 19
rect 1 -1 4 19
rect 10 -1 13 19
rect 19 -1 22 19
rect 28 -1 31 19
rect 37 -1 40 19
rect 61 -1 64 19
rect 78 -1 81 19
rect 87 -1 90 19
rect 104 -1 107 19
rect 113 -1 116 19
rect 130 -1 133 19
rect 139 -1 142 19
rect -8 -42 -6 -36
rect 0 -42 2 -36
rect 16 -42 18 -36
rect 78 -42 80 -36
rect 89 -42 91 -36
rect 113 -42 115 -36
<< ndiffusion >>
rect -9 -17 -8 -13
rect -11 -23 -8 -17
rect -5 -23 1 -13
rect 4 -20 10 -13
rect 4 -23 5 -20
rect 9 -23 10 -20
rect 13 -23 19 -13
rect 22 -17 23 -13
rect 22 -23 27 -17
rect 33 -19 36 -13
rect 35 -23 36 -19
rect 39 -23 43 -13
rect 46 -17 47 -13
rect 46 -23 51 -17
rect 58 -19 61 -13
rect 60 -23 61 -19
rect 64 -17 65 -13
rect 64 -23 67 -17
rect 75 -19 78 -13
rect 77 -23 78 -19
rect 81 -23 87 -13
rect 90 -17 91 -13
rect 90 -23 93 -17
rect 101 -19 104 -13
rect 103 -23 104 -19
rect 107 -23 113 -13
rect 116 -17 117 -13
rect 116 -23 119 -17
rect 127 -19 130 -13
rect 129 -23 130 -19
rect 133 -23 139 -13
rect 142 -17 143 -13
rect 142 -23 145 -17
rect 5 -73 8 -71
rect 7 -77 8 -73
rect 5 -95 8 -77
rect 10 -73 13 -71
rect 10 -77 11 -73
rect 10 -95 13 -77
rect 80 -83 83 -65
rect 82 -87 83 -83
rect 80 -89 83 -87
rect 85 -83 88 -65
rect 85 -87 86 -83
rect 85 -89 88 -87
<< pdiffusion >>
rect -11 17 -8 19
rect -9 9 -8 17
rect -11 -1 -8 9
rect -5 5 1 19
rect -5 1 -4 5
rect 0 1 1 5
rect -5 -1 1 1
rect 4 17 10 19
rect 4 9 5 17
rect 9 9 10 17
rect 4 -1 10 9
rect 13 5 19 19
rect 13 1 14 5
rect 18 1 19 5
rect 13 -1 19 1
rect 22 17 28 19
rect 22 9 23 17
rect 27 9 28 17
rect 22 -1 28 9
rect 31 5 37 19
rect 31 1 32 5
rect 36 1 37 5
rect 31 -1 37 1
rect 40 17 61 19
rect 40 10 41 17
rect 59 10 61 17
rect 40 -1 61 10
rect 64 6 67 19
rect 75 18 78 19
rect 77 9 78 18
rect 64 0 65 6
rect 64 -1 67 0
rect 75 -1 78 9
rect 81 10 87 19
rect 81 1 82 10
rect 86 1 87 10
rect 81 -1 87 1
rect 90 13 91 19
rect 95 13 104 19
rect 90 -1 104 13
rect 107 4 113 19
rect 107 0 108 4
rect 112 0 113 4
rect 107 -1 113 0
rect 116 14 117 19
rect 121 14 130 19
rect 116 -1 130 14
rect 133 4 139 19
rect 133 0 134 4
rect 138 0 139 4
rect 133 -1 139 0
rect 142 14 143 19
rect 142 -1 145 14
rect -11 -37 -8 -36
rect -9 -41 -8 -37
rect -11 -42 -8 -41
rect -6 -38 0 -36
rect -6 -42 -5 -38
rect -1 -42 0 -38
rect 2 -38 7 -36
rect 13 -38 16 -36
rect 2 -42 3 -38
rect 15 -42 16 -38
rect 18 -38 21 -36
rect 75 -38 78 -36
rect 18 -42 19 -38
rect 77 -42 78 -38
rect 80 -38 89 -36
rect 80 -42 81 -38
rect 85 -42 89 -38
rect 91 -38 94 -36
rect 110 -38 113 -36
rect 91 -42 92 -38
rect 112 -42 113 -38
rect 115 -38 118 -36
rect 115 -42 116 -38
<< ndcontact >>
rect -13 -17 -9 -13
rect 5 -24 9 -20
rect 23 -17 27 -13
rect 31 -23 35 -19
rect 47 -17 51 -13
rect 56 -23 60 -19
rect 65 -17 69 -13
rect 73 -23 77 -19
rect 91 -17 95 -13
rect 99 -23 103 -19
rect 117 -17 121 -13
rect 125 -23 129 -19
rect 143 -17 147 -13
rect 3 -77 7 -73
rect 11 -77 15 -73
rect 78 -87 82 -83
rect 86 -87 90 -83
<< pdcontact >>
rect -13 9 -9 17
rect -4 1 0 5
rect 5 9 9 17
rect 14 1 18 5
rect 23 9 27 17
rect 32 1 36 5
rect 41 10 59 17
rect 73 9 77 18
rect 65 0 69 6
rect 82 1 86 10
rect 91 13 95 19
rect 108 0 112 4
rect 117 14 121 19
rect 134 0 138 4
rect 143 14 147 19
rect -13 -41 -9 -37
rect -5 -42 -1 -38
rect 3 -42 7 -38
rect 11 -42 15 -38
rect 19 -42 23 -38
rect 73 -42 77 -38
rect 81 -42 85 -38
rect 92 -42 96 -38
rect 108 -42 112 -38
rect 116 -42 120 -38
<< psubstratepdiff >>
rect 78 -98 82 -94
<< nsubstratendiff >>
rect 211 35 220 44
<< polysilicon >>
rect -13 28 64 30
rect -8 19 -5 28
rect 1 19 4 20
rect 10 19 13 28
rect 19 19 22 20
rect 28 19 31 21
rect 37 19 40 21
rect 61 19 64 28
rect 78 19 81 21
rect 87 19 90 23
rect 104 19 107 21
rect 113 19 116 24
rect 130 19 133 21
rect 139 19 142 21
rect -8 -13 -5 -1
rect 1 -13 4 -1
rect 10 -13 13 -1
rect 19 -13 22 -1
rect 28 -8 31 -1
rect 37 -2 40 -1
rect 37 -4 47 -2
rect 43 -6 47 -4
rect 28 -12 35 -8
rect 36 -13 39 -12
rect 43 -13 46 -10
rect 61 -13 64 -1
rect 78 -2 81 -1
rect 80 -6 81 -2
rect 78 -13 81 -6
rect 87 -13 90 -1
rect 104 -3 107 -1
rect 104 -13 107 -7
rect 113 -13 116 -1
rect 130 -2 133 -1
rect 131 -6 133 -2
rect 130 -13 133 -6
rect 139 -2 142 -1
rect 139 -6 141 -2
rect 139 -13 142 -6
rect -8 -25 -5 -23
rect 1 -25 4 -23
rect 10 -25 13 -23
rect 19 -25 22 -23
rect 36 -25 39 -23
rect 43 -25 46 -23
rect 61 -25 64 -23
rect 78 -29 81 -23
rect 87 -25 90 -23
rect 104 -25 107 -23
rect 113 -25 116 -23
rect 130 -25 133 -23
rect 139 -25 142 -23
rect -8 -36 -6 -33
rect 0 -36 2 -33
rect 16 -36 18 -33
rect 78 -36 80 -33
rect 89 -36 91 -33
rect 113 -36 115 -33
rect -8 -44 -6 -42
rect 0 -44 2 -42
rect 16 -44 18 -42
rect 78 -44 80 -42
rect 89 -44 91 -42
rect 113 -44 115 -42
rect 83 -65 85 -64
rect 8 -71 10 -70
rect 83 -91 85 -89
rect 8 -97 10 -95
rect -297 -105 -294 -101
rect -290 -105 3 -101
rect 7 -105 53 -101
rect 57 -105 62 -101
rect -297 -461 62 -105
rect 65 -105 78 -101
rect 82 -105 121 -101
rect 125 -105 424 -101
rect 65 -461 424 -105
<< polycontact >>
rect -17 28 -13 32
rect 0 20 4 24
rect 19 20 23 24
rect 86 23 90 27
rect 112 24 116 28
rect 35 -12 39 -8
rect 43 -10 47 -6
rect 76 -6 80 -2
rect 103 -7 107 -3
rect 127 -6 131 -2
rect 141 -6 145 -2
rect -9 -33 -5 -29
rect -1 -33 3 -29
rect 15 -33 19 -29
rect 77 -33 81 -29
rect 88 -33 92 -29
rect 112 -33 116 -29
rect 82 -64 86 -60
rect 7 -70 11 -66
rect -294 -105 -290 -101
rect 3 -105 7 -101
rect 53 -105 57 -101
rect 78 -105 82 -101
rect 121 -105 125 -101
<< metal1 >>
rect 144 43 429 44
rect -299 35 -39 43
rect -33 35 429 43
rect -299 28 -17 32
rect 0 27 90 31
rect 0 24 4 27
rect -299 20 0 24
rect 89 19 147 20
rect 89 18 91 19
rect 30 17 73 18
rect -9 9 5 17
rect 9 9 23 17
rect 27 10 41 17
rect 59 10 73 17
rect 27 9 73 10
rect 77 13 91 18
rect 95 14 117 19
rect 121 14 143 19
rect 95 13 97 14
rect 77 9 79 13
rect 100 10 145 11
rect -13 1 -4 5
rect 18 1 27 5
rect 36 1 53 5
rect -13 -2 -9 1
rect -13 -13 -9 -6
rect 23 -8 27 1
rect 23 -12 35 -8
rect 23 -13 27 -12
rect 50 -13 53 1
rect -9 -29 -5 -13
rect -1 -17 23 -13
rect 51 -17 53 -13
rect 86 7 145 10
rect 86 6 105 7
rect 65 -2 69 0
rect 65 -6 72 -2
rect 83 -3 86 1
rect 112 0 121 4
rect 117 -2 121 0
rect 65 -13 69 -6
rect 83 -7 94 -3
rect 91 -9 94 -7
rect 117 -6 127 -2
rect 117 -13 121 -6
rect 134 -13 138 0
rect 141 -2 145 7
rect 134 -17 143 -13
rect -1 -29 2 -17
rect 9 -23 31 -20
rect 35 -23 56 -20
rect 60 -23 73 -20
rect 77 -23 99 -20
rect 103 -21 125 -20
rect 103 -23 121 -21
rect 134 -29 138 -17
rect 116 -33 138 -29
rect -13 -59 -9 -41
rect 3 -52 7 -42
rect 23 -42 61 -38
rect 3 -56 21 -52
rect 40 -59 44 -49
rect 57 -53 61 -42
rect 81 -45 85 -42
rect 108 -45 112 -42
rect 81 -49 105 -45
rect 109 -49 112 -45
rect 116 -53 120 -42
rect 57 -57 120 -53
rect -13 -63 44 -59
rect 15 -67 19 -63
rect 15 -71 426 -67
rect 3 -101 7 -77
rect -302 -105 -294 -101
rect 15 -77 19 -71
rect 11 -113 15 -77
rect 33 -78 105 -74
rect 78 -101 82 -87
rect 57 -105 78 -101
rect 94 -87 426 -83
rect 86 -111 90 -87
rect 121 -101 125 -96
<< m2contact >>
rect -39 35 -33 43
rect 23 20 27 24
rect 108 24 112 28
rect -17 9 -13 17
rect -13 -6 -9 -2
rect 43 -6 47 -2
rect 43 -17 47 -13
rect 72 -6 76 -2
rect 91 -13 95 -9
rect 103 -11 107 -7
rect 121 -25 125 -21
rect 19 -33 23 -29
rect 81 -33 85 -29
rect 92 -33 96 -29
rect -5 -46 -1 -42
rect 69 -42 73 -38
rect 96 -42 100 -38
rect 11 -46 15 -42
rect 40 -49 44 -45
rect 21 -56 25 -52
rect 105 -49 109 -45
rect 3 -70 7 -66
rect 78 -64 82 -60
rect 29 -78 33 -74
rect 105 -78 109 -74
rect 90 -87 94 -83
rect 121 -96 125 -92
<< metal2 >>
rect -39 17 -33 35
rect 12 20 23 24
rect 27 20 112 24
rect -39 9 -17 17
rect 12 6 16 20
rect -298 2 17 6
rect -9 -6 43 -2
rect 76 -3 103 -2
rect 76 -6 107 -3
rect 98 -7 107 -6
rect 81 -13 91 -9
rect 43 -29 47 -17
rect 23 -33 47 -29
rect 81 -29 85 -13
rect 103 -23 107 -11
rect 92 -27 107 -23
rect 92 -29 96 -27
rect 63 -42 69 -38
rect -297 -46 -5 -45
rect -1 -46 11 -45
rect 63 -45 67 -42
rect -297 -49 15 -46
rect 44 -49 67 -45
rect 96 -52 100 -42
rect 25 -56 100 -52
rect -298 -63 33 -59
rect -297 -70 3 -66
rect 29 -74 33 -63
rect 61 -64 78 -60
rect 61 -81 65 -64
rect -297 -85 65 -81
rect 90 -83 94 -56
rect 105 -74 109 -49
rect 121 -92 125 -25
<< labels >>
rlabel metal1 -4 15 -4 15 1 Vdd
rlabel polycontact 2 20 3 21 1 C1?
rlabel polycontact 20 20 21 21 1 C2?
rlabel metal1 28 -22 28 -22 1 Gnd
rlabel metal1 95 -48 95 -48 1 Iref
rlabel metal2 -2 -48 -2 -48 1 Iin
rlabel metal2 -29 -69 -29 -69 1 CLC1
rlabel metal2 92 -79 92 -79 1 VC2
rlabel metal1 13 -98 13 -98 1 VC1
rlabel metal1 4 -99 4 -99 1 Gnd
rlabel polysilicon -7 29 -7 29 1 Iin?
rlabel metal2 -35 3 -35 3 1 C2?
rlabel metal2 -29 -84 -29 -84 1 CLC2
rlabel metal2 -294 -61 -294 -61 1 Iref
<< end >>
