magic
tech scmos
timestamp 1355680695
<< nwell >>
rect -1243 3082 -1239 3103
<< pwell >>
rect -868 2952 -864 2963
rect -1067 2931 -997 2936
<< metal1 >>
rect -193 3184 379 3195
rect -977 3111 -905 3121
rect -1243 3082 -1239 3099
rect -1029 3097 -1019 3101
rect -978 3097 -949 3101
rect -1029 3076 -1025 3097
rect -914 3076 -905 3111
rect -193 3095 -183 3184
rect -914 3072 -909 3076
rect 128 3039 144 3056
rect 128 3001 151 3039
rect -135 2903 -100 2918
rect 196 2740 209 3123
rect 369 3107 379 3184
rect 357 3086 379 3107
rect 196 2726 197 2740
rect 226 2690 242 2894
rect 164 2661 200 2665
rect -787 2604 3 2619
rect 169 2592 222 2597
rect -101 2571 328 2575
rect 336 2514 360 2582
rect 377 2575 381 2582
rect 374 2571 381 2575
rect 377 2522 381 2571
rect 386 2531 391 2581
rect 386 2525 463 2531
rect 377 2517 436 2522
rect -874 2188 -843 2230
rect -8 1597 10 2507
rect 336 2494 410 2514
rect 177 1953 185 2133
rect 300 1611 301 1622
rect 305 1611 306 1622
rect 259 1563 274 1611
rect 300 1607 306 1611
rect 300 1563 306 1566
rect 325 1564 348 1611
rect 300 1552 301 1563
rect 305 1552 306 1563
rect 392 1529 400 1684
rect 418 1622 436 2517
rect 423 1611 436 1622
rect 418 1563 436 1611
rect 406 1554 436 1563
rect 406 1529 414 1554
rect -12 1507 4 1512
rect 445 1511 463 2525
rect -2597 1005 -2585 1021
rect 19 -9 37 19
rect 48 0 79 7
rect 48 -8 52 0
rect 129 -7 152 16
rect 65 -17 152 -7
rect 47 -75 51 -52
<< m2contact >>
rect -1243 3099 -1239 3103
rect -1029 3072 -1025 3076
rect 196 3123 209 3142
rect -909 3072 -905 3076
rect -81 3039 -74 3056
rect 144 3039 151 3056
rect -868 2952 -864 2963
rect -100 2903 -95 2918
rect 14 2904 18 2918
rect 197 2726 209 2740
rect 159 2661 164 2665
rect 238 2661 243 2665
rect -798 2604 -787 2619
rect 3 2603 9 2619
rect 222 2590 230 2597
rect 18 2580 45 2587
rect -107 2571 -101 2575
rect 328 2571 332 2575
rect 368 2580 373 2584
rect 370 2571 374 2575
rect 19 2504 46 2511
rect 70 2482 87 2494
rect 177 2133 185 2140
rect 382 1684 400 1701
rect 301 1611 305 1622
rect 301 1552 305 1563
rect -13 1521 -8 1540
rect 19 1521 24 1540
rect 418 1611 423 1622
rect -56 1507 -51 1512
rect 177 1501 185 1511
rect 445 1499 463 1511
rect -12 1487 -8 1494
rect 146 1487 152 1494
<< metal2 >>
rect -1253 3089 -1246 3128
rect -1243 3123 196 3142
rect -1243 3103 -1236 3123
rect -1239 3099 -1236 3103
rect -1025 3072 -987 3076
rect -992 3006 -987 3072
rect -909 3069 -905 3072
rect -909 3065 -864 3069
rect -1001 3001 -987 3006
rect -1001 2936 -997 3001
rect -868 2963 -864 3065
rect -74 3039 144 3056
rect -1067 2931 -997 2936
rect -95 2904 14 2918
rect -95 2903 8 2904
rect 180 2740 209 2741
rect 180 2726 197 2740
rect 179 2661 238 2665
rect -392 2495 -386 2625
rect -107 2575 -101 2625
rect 3 2619 9 2628
rect 18 2511 45 2580
rect 18 2504 19 2511
rect 158 2509 164 2581
rect 179 2514 184 2582
rect 171 2509 184 2514
rect -392 2494 87 2495
rect -392 2482 70 2494
rect 222 2140 230 2590
rect 373 2580 385 2584
rect 332 2571 370 2575
rect 381 2517 385 2580
rect 185 2133 230 2140
rect 368 1701 385 2517
rect 368 1684 382 1701
rect 305 1611 418 1622
rect 305 1552 386 1563
rect -8 1521 19 1540
rect 378 1512 386 1552
rect -51 1511 185 1512
rect -51 1507 177 1511
rect -56 1502 177 1507
rect 378 1511 463 1512
rect 378 1499 445 1511
rect -8 1487 146 1494
use NOT  NOT_4
timestamp 1355475633
transform -1 0 -978 0 -1 3107
box -5 -23 43 41
use stateMachine  stateMachine_0
timestamp 1355540337
transform 1 0 -1265 0 1 3050
box -14 -441 1196 68
use NOT  NOT_3
timestamp 1355475633
transform -1 0 238 0 -1 2671
box -5 -23 43 41
use msb_registers  msb_registers_0
timestamp 1355455137
transform 0 1 227 1 0 2875
box -295 -224 301 222
use Comparator  Comparator_0
timestamp 1355605154
transform 0 1 -1060 1 0 1639
box -6 -28 815 195
use AnalogSwitch  AnalogSwitch_0
timestamp 1355620377
transform 0 1 -256 -1 0 2054
box -325 -461 424 47
use NOT  NOT_2
timestamp 1355475633
transform 0 1 295 -1 0 1606
box -5 -23 43 41
use NOT  NOT_1
timestamp 1355475633
transform -1 0 -13 0 -1 1517
box -5 -23 43 41
use lsb_registers_Layout  lsb_registers_Layout_0
timestamp 1355674588
transform 0 1 263 -1 0 1521
box -990 -263 1521 160
use NOT  NOT_0
timestamp 1355475633
transform 0 1 42 -1 0 -12
box -5 -23 43 41
<< labels >>
rlabel metal1 49 -72 49 -72 1 GO?
rlabel metal2 -1250 3125 -1250 3125 1 CO
rlabel metal2 -1240 3124 -1240 3124 1 CLK
<< end >>
