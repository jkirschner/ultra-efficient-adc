magic
tech scmos
timestamp 1354990610
<< nwell >>
rect 213 -299 316 -208
rect 322 -274 425 -208
<< pwell >>
rect 213 -344 316 -299
rect 322 -344 425 -274
<< ntransistor >>
rect 335 -295 338 -285
rect 342 -295 345 -285
rect 351 -295 354 -285
rect 358 -295 361 -285
rect 367 -295 370 -285
rect 374 -295 377 -285
rect 383 -295 386 -285
rect 390 -295 393 -285
rect 399 -291 402 -281
rect 226 -320 229 -310
rect 233 -320 236 -310
rect 242 -320 245 -310
rect 249 -320 252 -310
rect 258 -320 261 -310
rect 265 -320 268 -310
rect 274 -320 277 -310
rect 281 -320 284 -310
rect 290 -316 293 -306
rect 352 -308 362 -305
rect 382 -308 392 -305
rect 402 -308 405 -298
rect 243 -333 253 -330
rect 273 -333 283 -330
rect 293 -333 296 -323
rect 337 -333 340 -318
rect 346 -333 349 -318
rect 355 -333 358 -318
rect 364 -333 367 -318
rect 373 -333 376 -318
rect 382 -333 385 -318
rect 391 -333 394 -318
rect 400 -333 403 -318
<< ptransistor >>
rect 224 -262 227 -220
rect 233 -246 236 -220
rect 242 -246 245 -220
rect 251 -246 254 -220
rect 236 -258 256 -255
rect 263 -262 266 -220
rect 272 -246 275 -220
rect 281 -246 284 -220
rect 290 -246 293 -220
rect 345 -233 365 -230
rect 384 -233 404 -230
rect 275 -258 295 -255
rect 226 -289 229 -269
rect 233 -289 236 -269
rect 242 -289 245 -269
rect 249 -289 252 -269
rect 258 -289 261 -269
rect 265 -289 268 -269
rect 274 -289 277 -269
rect 281 -289 284 -269
rect 290 -293 293 -273
rect 302 -282 305 -262
rect 335 -264 338 -244
rect 342 -264 345 -244
rect 351 -264 354 -244
rect 358 -264 361 -244
rect 367 -264 370 -244
rect 374 -264 377 -244
rect 383 -264 386 -244
rect 390 -264 393 -244
rect 399 -268 402 -248
rect 411 -257 414 -237
<< ndiffusion >>
rect 396 -285 399 -281
rect 330 -286 335 -285
rect 334 -294 335 -286
rect 330 -295 335 -294
rect 338 -295 342 -285
rect 345 -290 351 -285
rect 345 -294 346 -290
rect 350 -294 351 -290
rect 345 -295 351 -294
rect 354 -295 358 -285
rect 361 -286 367 -285
rect 361 -294 362 -286
rect 366 -294 367 -286
rect 361 -295 367 -294
rect 370 -295 374 -285
rect 377 -290 383 -285
rect 377 -294 378 -290
rect 382 -294 383 -290
rect 377 -295 383 -294
rect 386 -295 390 -285
rect 393 -286 399 -285
rect 393 -294 394 -286
rect 398 -291 399 -286
rect 402 -282 408 -281
rect 402 -286 403 -282
rect 407 -286 408 -282
rect 402 -291 408 -286
rect 393 -295 398 -294
rect 352 -304 353 -300
rect 357 -304 362 -300
rect 352 -305 362 -304
rect 399 -299 402 -298
rect 382 -304 383 -300
rect 391 -304 392 -300
rect 382 -305 392 -304
rect 287 -310 290 -306
rect 219 -311 226 -310
rect 219 -319 221 -311
rect 225 -319 226 -311
rect 219 -320 226 -319
rect 229 -320 233 -310
rect 236 -315 242 -310
rect 236 -319 237 -315
rect 241 -319 242 -315
rect 236 -320 242 -319
rect 245 -320 249 -310
rect 252 -311 258 -310
rect 252 -319 253 -311
rect 257 -319 258 -311
rect 252 -320 258 -319
rect 261 -320 265 -310
rect 268 -315 274 -310
rect 268 -319 269 -315
rect 273 -319 274 -315
rect 268 -320 274 -319
rect 277 -320 281 -310
rect 284 -311 290 -310
rect 284 -319 285 -311
rect 289 -316 290 -311
rect 293 -307 299 -306
rect 293 -311 294 -307
rect 298 -311 299 -307
rect 401 -307 402 -299
rect 399 -308 402 -307
rect 405 -300 409 -298
rect 405 -307 406 -300
rect 405 -308 409 -307
rect 293 -316 299 -311
rect 352 -309 362 -308
rect 352 -313 353 -309
rect 361 -313 362 -309
rect 382 -309 392 -308
rect 382 -313 383 -309
rect 391 -313 392 -309
rect 284 -320 289 -319
rect 243 -329 244 -325
rect 248 -329 253 -325
rect 243 -330 253 -329
rect 332 -322 337 -318
rect 290 -324 293 -323
rect 273 -329 274 -325
rect 282 -329 283 -325
rect 273 -330 283 -329
rect 292 -332 293 -324
rect 290 -333 293 -332
rect 296 -325 300 -323
rect 296 -332 297 -325
rect 336 -326 337 -322
rect 332 -328 337 -326
rect 336 -332 337 -328
rect 296 -333 300 -332
rect 332 -333 337 -332
rect 340 -319 346 -318
rect 340 -323 341 -319
rect 345 -323 346 -319
rect 340 -333 346 -323
rect 349 -326 355 -318
rect 349 -332 350 -326
rect 354 -332 355 -326
rect 349 -333 355 -332
rect 358 -319 364 -318
rect 358 -323 359 -319
rect 363 -323 364 -319
rect 358 -333 364 -323
rect 367 -319 373 -318
rect 367 -332 368 -319
rect 372 -332 373 -319
rect 367 -333 373 -332
rect 376 -319 382 -318
rect 376 -323 377 -319
rect 381 -323 382 -319
rect 376 -333 382 -323
rect 385 -326 391 -318
rect 385 -332 386 -326
rect 390 -332 391 -326
rect 385 -333 391 -332
rect 394 -319 400 -318
rect 394 -323 395 -319
rect 399 -323 400 -319
rect 394 -333 400 -323
rect 403 -322 408 -318
rect 403 -326 404 -322
rect 403 -328 408 -326
rect 403 -332 404 -328
rect 403 -333 408 -332
rect 243 -334 253 -333
rect 243 -338 244 -334
rect 252 -338 253 -334
rect 273 -334 283 -333
rect 273 -338 274 -334
rect 282 -338 283 -334
<< pdiffusion >>
rect 219 -227 224 -220
rect 223 -231 224 -227
rect 219 -241 224 -231
rect 223 -245 224 -241
rect 221 -262 224 -245
rect 227 -221 233 -220
rect 227 -225 228 -221
rect 232 -225 233 -221
rect 227 -234 233 -225
rect 227 -238 228 -234
rect 232 -238 233 -234
rect 227 -246 233 -238
rect 236 -227 242 -220
rect 236 -231 237 -227
rect 241 -231 242 -227
rect 236 -241 242 -231
rect 236 -245 237 -241
rect 241 -245 242 -241
rect 236 -246 242 -245
rect 245 -221 251 -220
rect 245 -225 246 -221
rect 250 -225 251 -221
rect 245 -234 251 -225
rect 245 -238 246 -234
rect 250 -238 251 -234
rect 245 -246 251 -238
rect 254 -227 263 -220
rect 254 -231 255 -227
rect 262 -231 263 -227
rect 254 -241 263 -231
rect 254 -245 255 -241
rect 262 -245 263 -241
rect 254 -246 263 -245
rect 227 -250 231 -246
rect 227 -254 228 -250
rect 236 -254 237 -250
rect 227 -262 230 -254
rect 236 -255 256 -254
rect 236 -259 256 -258
rect 236 -261 240 -259
rect 247 -261 256 -259
rect 260 -262 263 -246
rect 266 -221 272 -220
rect 266 -225 267 -221
rect 271 -225 272 -221
rect 266 -234 272 -225
rect 266 -238 267 -234
rect 271 -238 272 -234
rect 266 -246 272 -238
rect 275 -227 281 -220
rect 275 -231 276 -227
rect 280 -231 281 -227
rect 275 -241 281 -231
rect 275 -245 276 -241
rect 280 -245 281 -241
rect 275 -246 281 -245
rect 284 -221 290 -220
rect 284 -225 285 -221
rect 289 -225 290 -221
rect 284 -234 290 -225
rect 284 -238 285 -234
rect 289 -238 290 -234
rect 284 -246 290 -238
rect 293 -227 297 -220
rect 293 -231 294 -227
rect 345 -229 346 -225
rect 345 -230 365 -229
rect 384 -229 385 -225
rect 384 -230 404 -229
rect 293 -241 297 -231
rect 345 -234 365 -233
rect 345 -236 349 -234
rect 356 -236 365 -234
rect 384 -234 404 -233
rect 384 -236 386 -234
rect 390 -236 404 -234
rect 293 -245 294 -241
rect 408 -240 411 -237
rect 410 -244 411 -240
rect 328 -245 335 -244
rect 293 -246 297 -245
rect 266 -250 270 -246
rect 266 -254 267 -250
rect 275 -254 276 -250
rect 266 -262 269 -254
rect 275 -255 295 -254
rect 328 -254 330 -245
rect 334 -254 335 -245
rect 328 -256 335 -254
rect 275 -259 295 -258
rect 275 -261 277 -259
rect 281 -261 295 -259
rect 299 -265 302 -262
rect 301 -269 302 -265
rect 219 -270 226 -269
rect 219 -279 221 -270
rect 225 -279 226 -270
rect 219 -281 226 -279
rect 223 -289 226 -281
rect 229 -289 233 -269
rect 236 -271 242 -269
rect 236 -277 237 -271
rect 241 -277 242 -271
rect 236 -281 242 -277
rect 236 -287 237 -281
rect 241 -287 242 -281
rect 236 -289 242 -287
rect 245 -289 249 -269
rect 252 -271 258 -269
rect 252 -288 253 -271
rect 257 -288 258 -271
rect 252 -289 258 -288
rect 261 -289 265 -269
rect 268 -271 274 -269
rect 268 -277 269 -271
rect 273 -277 274 -271
rect 268 -281 274 -277
rect 268 -287 269 -281
rect 273 -287 274 -281
rect 268 -289 274 -287
rect 277 -289 281 -269
rect 284 -271 289 -269
rect 284 -287 285 -271
rect 289 -287 290 -273
rect 284 -289 290 -287
rect 287 -293 290 -289
rect 293 -286 296 -273
rect 299 -282 302 -269
rect 305 -263 308 -262
rect 305 -281 306 -263
rect 332 -264 335 -256
rect 338 -264 342 -244
rect 345 -246 351 -244
rect 345 -252 346 -246
rect 350 -252 351 -246
rect 345 -256 351 -252
rect 345 -262 346 -256
rect 350 -262 351 -256
rect 345 -264 351 -262
rect 354 -264 358 -244
rect 361 -246 367 -244
rect 361 -263 362 -246
rect 366 -263 367 -246
rect 361 -264 367 -263
rect 370 -264 374 -244
rect 377 -246 383 -244
rect 377 -252 378 -246
rect 382 -252 383 -246
rect 377 -256 383 -252
rect 377 -262 378 -256
rect 382 -262 383 -256
rect 377 -264 383 -262
rect 386 -264 390 -244
rect 393 -246 398 -244
rect 393 -262 394 -246
rect 398 -262 399 -248
rect 393 -264 399 -262
rect 305 -282 308 -281
rect 396 -268 399 -264
rect 402 -261 405 -248
rect 408 -257 411 -244
rect 414 -238 417 -237
rect 414 -256 415 -238
rect 414 -257 417 -256
rect 402 -262 408 -261
rect 402 -266 403 -262
rect 407 -266 408 -262
rect 402 -268 408 -266
rect 293 -287 299 -286
rect 293 -291 294 -287
rect 298 -291 299 -287
rect 293 -293 299 -291
<< ndcontact >>
rect 330 -294 334 -286
rect 346 -294 350 -290
rect 362 -294 366 -286
rect 378 -294 382 -290
rect 394 -294 398 -286
rect 403 -286 407 -282
rect 353 -304 357 -300
rect 383 -304 391 -300
rect 221 -319 225 -311
rect 237 -319 241 -315
rect 253 -319 257 -311
rect 269 -319 273 -315
rect 285 -319 289 -311
rect 294 -311 298 -307
rect 397 -307 401 -299
rect 406 -307 410 -300
rect 353 -313 361 -309
rect 383 -313 391 -309
rect 244 -329 248 -325
rect 274 -329 282 -325
rect 288 -332 292 -324
rect 297 -332 301 -325
rect 332 -326 336 -322
rect 332 -332 336 -328
rect 341 -323 345 -319
rect 350 -332 354 -326
rect 359 -323 363 -319
rect 368 -332 372 -319
rect 377 -323 381 -319
rect 386 -332 390 -326
rect 395 -323 399 -319
rect 404 -326 408 -322
rect 404 -332 408 -328
rect 244 -338 252 -334
rect 274 -338 282 -334
<< pdcontact >>
rect 219 -231 223 -227
rect 219 -245 223 -241
rect 228 -225 232 -221
rect 228 -238 232 -234
rect 237 -231 241 -227
rect 237 -245 241 -241
rect 246 -225 250 -221
rect 246 -238 250 -234
rect 255 -231 262 -227
rect 255 -245 262 -241
rect 228 -254 232 -250
rect 237 -254 256 -250
rect 240 -263 247 -259
rect 267 -225 271 -221
rect 267 -238 271 -234
rect 276 -231 280 -227
rect 276 -245 280 -241
rect 285 -225 289 -221
rect 285 -238 289 -234
rect 294 -231 298 -227
rect 346 -229 365 -225
rect 385 -229 404 -225
rect 349 -238 356 -234
rect 386 -238 390 -234
rect 294 -245 298 -241
rect 406 -244 410 -240
rect 267 -254 271 -250
rect 276 -254 295 -250
rect 330 -254 334 -245
rect 277 -263 281 -259
rect 297 -269 301 -265
rect 221 -279 225 -270
rect 237 -277 241 -271
rect 237 -287 241 -281
rect 253 -288 257 -271
rect 269 -277 273 -271
rect 269 -287 273 -281
rect 285 -287 289 -271
rect 306 -281 310 -263
rect 346 -252 350 -246
rect 346 -262 350 -256
rect 362 -263 366 -246
rect 378 -252 382 -246
rect 378 -262 382 -256
rect 394 -262 398 -246
rect 415 -256 419 -238
rect 403 -266 407 -262
rect 294 -291 298 -287
<< psubstratepdiff >>
rect 222 -336 226 -332
<< nsubstratendiff >>
rect 307 -221 311 -217
rect 416 -222 420 -218
<< psubstratepcontact >>
rect 226 -336 230 -332
<< nsubstratencontact >>
rect 303 -221 307 -217
rect 412 -222 416 -218
<< polysilicon >>
rect 224 -218 228 -216
rect 232 -218 237 -216
rect 241 -218 246 -216
rect 250 -218 267 -216
rect 271 -218 276 -216
rect 280 -218 285 -216
rect 289 -218 293 -216
rect 224 -219 293 -218
rect 224 -220 227 -219
rect 233 -220 236 -219
rect 242 -220 245 -219
rect 251 -220 254 -219
rect 263 -220 266 -219
rect 272 -220 275 -219
rect 281 -220 284 -219
rect 290 -220 293 -219
rect 233 -248 236 -246
rect 242 -248 245 -246
rect 251 -248 254 -246
rect 231 -258 236 -255
rect 256 -258 258 -255
rect 224 -264 227 -262
rect 340 -233 345 -230
rect 365 -233 367 -230
rect 380 -233 384 -230
rect 404 -233 414 -230
rect 411 -237 414 -233
rect 335 -244 338 -242
rect 342 -244 345 -242
rect 351 -244 354 -242
rect 358 -244 361 -242
rect 367 -244 370 -242
rect 374 -244 377 -242
rect 383 -244 386 -242
rect 390 -244 393 -239
rect 272 -248 275 -246
rect 281 -248 284 -246
rect 290 -248 293 -246
rect 270 -258 275 -255
rect 295 -258 305 -255
rect 263 -264 266 -262
rect 302 -262 305 -258
rect 226 -269 229 -267
rect 233 -269 236 -267
rect 242 -269 245 -267
rect 249 -269 252 -267
rect 258 -269 261 -267
rect 265 -269 268 -267
rect 274 -269 277 -267
rect 281 -269 284 -264
rect 290 -273 293 -271
rect 226 -297 229 -289
rect 233 -304 236 -289
rect 242 -291 245 -289
rect 249 -291 252 -289
rect 226 -310 229 -308
rect 233 -310 236 -308
rect 242 -310 245 -295
rect 258 -298 261 -289
rect 265 -291 268 -289
rect 249 -310 252 -302
rect 258 -310 261 -308
rect 265 -310 268 -295
rect 274 -304 277 -289
rect 281 -291 284 -289
rect 399 -248 402 -246
rect 335 -272 338 -264
rect 342 -279 345 -264
rect 351 -266 354 -264
rect 358 -266 361 -264
rect 302 -284 305 -282
rect 335 -285 338 -283
rect 342 -285 345 -283
rect 351 -285 354 -270
rect 367 -273 370 -264
rect 374 -266 377 -264
rect 358 -285 361 -277
rect 367 -285 370 -283
rect 374 -285 377 -270
rect 383 -279 386 -264
rect 390 -266 393 -264
rect 411 -259 414 -257
rect 399 -269 402 -268
rect 383 -285 386 -283
rect 390 -285 393 -277
rect 399 -281 402 -273
rect 290 -294 293 -293
rect 399 -293 402 -291
rect 335 -297 338 -295
rect 342 -297 345 -295
rect 351 -297 354 -295
rect 358 -297 361 -295
rect 274 -310 277 -308
rect 281 -310 284 -302
rect 290 -306 293 -298
rect 334 -301 338 -297
rect 367 -301 370 -295
rect 374 -297 377 -295
rect 383 -297 386 -295
rect 390 -297 393 -295
rect 402 -298 405 -296
rect 367 -305 368 -301
rect 346 -308 352 -305
rect 362 -308 364 -305
rect 376 -308 382 -305
rect 392 -308 396 -305
rect 393 -309 396 -308
rect 402 -309 405 -308
rect 393 -312 405 -309
rect 290 -318 293 -316
rect 337 -318 340 -316
rect 346 -318 349 -316
rect 355 -318 358 -316
rect 364 -318 367 -316
rect 373 -318 376 -316
rect 382 -318 385 -316
rect 391 -318 394 -316
rect 400 -318 403 -316
rect 226 -322 229 -320
rect 233 -322 236 -320
rect 242 -322 245 -320
rect 249 -322 252 -320
rect 258 -326 261 -320
rect 265 -322 268 -320
rect 274 -322 277 -320
rect 281 -322 284 -320
rect 293 -323 296 -321
rect 258 -330 259 -326
rect 237 -333 243 -330
rect 253 -333 255 -330
rect 267 -333 273 -330
rect 283 -333 287 -330
rect 284 -334 287 -333
rect 293 -334 296 -333
rect 284 -337 296 -334
rect 337 -334 340 -333
rect 346 -334 349 -333
rect 355 -334 358 -333
rect 364 -334 367 -333
rect 373 -334 376 -333
rect 382 -334 385 -333
rect 391 -334 394 -333
rect 400 -334 403 -333
rect 337 -337 403 -334
rect 337 -339 341 -337
rect 345 -339 350 -337
rect 354 -339 359 -337
rect 363 -339 377 -337
rect 381 -339 386 -337
rect 390 -339 395 -337
rect 399 -339 403 -337
<< polycontact >>
rect 228 -218 232 -214
rect 237 -218 241 -214
rect 246 -218 250 -214
rect 267 -218 271 -214
rect 276 -218 280 -214
rect 285 -218 289 -214
rect 231 -262 235 -258
rect 340 -237 344 -233
rect 379 -237 383 -233
rect 358 -242 362 -238
rect 393 -242 397 -238
rect 270 -262 274 -258
rect 249 -267 253 -263
rect 284 -267 288 -263
rect 225 -301 229 -297
rect 241 -295 245 -291
rect 233 -308 237 -304
rect 249 -302 253 -298
rect 257 -302 261 -298
rect 265 -295 269 -291
rect 334 -276 338 -272
rect 350 -270 354 -266
rect 342 -283 346 -279
rect 358 -277 362 -273
rect 366 -277 370 -273
rect 374 -270 378 -266
rect 399 -273 403 -269
rect 382 -283 386 -279
rect 390 -277 394 -273
rect 290 -298 294 -294
rect 273 -308 277 -304
rect 281 -302 285 -298
rect 330 -301 334 -297
rect 346 -305 350 -301
rect 368 -305 372 -301
rect 376 -305 380 -301
rect 225 -326 229 -322
rect 237 -330 241 -326
rect 259 -330 263 -326
rect 267 -330 271 -326
rect 341 -341 345 -337
rect 350 -341 354 -337
rect 359 -341 363 -337
rect 377 -341 381 -337
rect 386 -341 390 -337
rect 395 -341 399 -337
<< metal1 >>
rect 213 -227 223 -211
rect 242 -213 246 -208
rect 228 -214 289 -213
rect 232 -216 237 -214
rect 241 -216 246 -214
rect 250 -216 267 -214
rect 271 -216 276 -214
rect 280 -216 285 -214
rect 294 -216 316 -211
rect 293 -217 316 -216
rect 293 -221 303 -217
rect 307 -221 316 -217
rect 232 -224 246 -221
rect 254 -227 263 -221
rect 271 -224 285 -221
rect 293 -227 316 -221
rect 213 -231 219 -227
rect 223 -231 237 -228
rect 254 -228 255 -227
rect 241 -231 255 -228
rect 262 -228 263 -227
rect 262 -231 276 -228
rect 293 -228 294 -227
rect 280 -231 294 -228
rect 298 -231 316 -227
rect 213 -234 224 -231
rect 217 -241 224 -234
rect 232 -238 246 -234
rect 254 -241 263 -231
rect 293 -234 316 -231
rect 322 -218 425 -211
rect 322 -222 412 -218
rect 416 -222 425 -218
rect 322 -225 425 -222
rect 322 -229 346 -225
rect 365 -229 385 -225
rect 404 -229 425 -225
rect 322 -234 334 -229
rect 271 -238 285 -234
rect 293 -241 307 -234
rect 217 -245 219 -241
rect 223 -245 237 -241
rect 241 -245 255 -241
rect 262 -245 276 -241
rect 280 -245 294 -241
rect 298 -245 307 -241
rect 217 -247 307 -245
rect 217 -256 225 -247
rect 236 -250 264 -247
rect 275 -250 307 -247
rect 215 -282 218 -259
rect 221 -270 225 -256
rect 236 -254 237 -250
rect 256 -254 264 -250
rect 275 -254 276 -250
rect 295 -254 307 -250
rect 330 -245 334 -234
rect 340 -246 344 -237
rect 356 -238 358 -234
rect 340 -250 346 -246
rect 228 -258 232 -254
rect 228 -262 231 -258
rect 228 -271 232 -262
rect 247 -263 249 -259
rect 228 -275 237 -271
rect 215 -297 221 -282
rect 257 -276 261 -254
rect 267 -258 271 -254
rect 267 -262 270 -258
rect 267 -271 272 -262
rect 281 -267 284 -263
rect 291 -265 295 -254
rect 306 -263 313 -262
rect 291 -269 297 -265
rect 291 -271 295 -269
rect 267 -273 269 -271
rect 289 -276 295 -271
rect 310 -285 313 -263
rect 324 -272 330 -262
rect 366 -251 370 -229
rect 378 -237 379 -233
rect 400 -234 425 -229
rect 378 -246 382 -237
rect 390 -242 393 -238
rect 400 -240 404 -234
rect 400 -244 406 -240
rect 400 -246 404 -244
rect 398 -251 404 -246
rect 415 -262 419 -260
rect 407 -266 411 -262
rect 354 -269 362 -266
rect 366 -269 374 -266
rect 324 -276 334 -272
rect 338 -276 358 -273
rect 324 -283 330 -276
rect 374 -276 390 -273
rect 346 -283 382 -280
rect 406 -282 411 -266
rect 415 -267 422 -262
rect 298 -288 300 -287
rect 298 -291 313 -288
rect 245 -294 253 -291
rect 257 -294 265 -291
rect 215 -301 225 -297
rect 229 -301 249 -298
rect 215 -308 221 -301
rect 265 -301 281 -298
rect 237 -308 273 -305
rect 297 -307 313 -291
rect 298 -311 313 -307
rect 324 -311 327 -283
rect 334 -294 343 -286
rect 337 -309 343 -294
rect 219 -317 221 -311
rect 213 -319 221 -317
rect 213 -329 222 -319
rect 237 -326 241 -319
rect 251 -319 253 -311
rect 213 -332 234 -329
rect 213 -336 226 -332
rect 230 -333 234 -332
rect 251 -333 255 -319
rect 267 -322 273 -319
rect 330 -316 343 -309
rect 346 -301 350 -294
rect 360 -294 362 -286
rect 330 -317 337 -316
rect 267 -326 271 -322
rect 285 -323 289 -319
rect 285 -324 290 -323
rect 285 -332 288 -324
rect 285 -333 290 -332
rect 230 -334 290 -333
rect 230 -336 244 -334
rect 213 -338 244 -336
rect 252 -338 274 -334
rect 282 -335 290 -334
rect 308 -335 316 -317
rect 282 -338 316 -335
rect 213 -344 316 -338
rect 322 -322 337 -317
rect 346 -319 349 -305
rect 360 -308 364 -294
rect 376 -297 382 -294
rect 407 -288 411 -282
rect 417 -285 422 -267
rect 407 -294 422 -288
rect 376 -301 380 -297
rect 394 -298 398 -294
rect 394 -299 399 -298
rect 353 -309 373 -308
rect 361 -313 373 -309
rect 367 -319 373 -313
rect 322 -326 332 -322
rect 336 -326 337 -322
rect 345 -323 359 -319
rect 367 -326 368 -319
rect 322 -328 350 -326
rect 322 -332 332 -328
rect 336 -332 350 -328
rect 354 -332 368 -326
rect 372 -326 373 -319
rect 376 -319 379 -305
rect 394 -307 397 -299
rect 394 -308 399 -307
rect 382 -309 399 -308
rect 382 -313 383 -309
rect 391 -310 399 -309
rect 391 -313 409 -310
rect 417 -311 422 -294
rect 382 -314 409 -313
rect 404 -317 409 -314
rect 376 -323 377 -319
rect 381 -323 395 -319
rect 404 -322 425 -317
rect 408 -326 425 -322
rect 372 -332 386 -326
rect 390 -328 425 -326
rect 390 -332 404 -328
rect 408 -332 425 -328
rect 322 -334 425 -332
rect 322 -344 336 -334
rect 345 -341 350 -339
rect 354 -341 359 -339
rect 363 -341 377 -339
rect 381 -341 386 -339
rect 390 -341 395 -339
rect 341 -342 399 -341
rect 355 -344 359 -342
rect 381 -344 385 -342
rect 404 -344 425 -334
<< m2contact >>
rect 353 -242 358 -238
rect 244 -267 249 -263
rect 237 -281 241 -277
rect 277 -267 281 -263
rect 346 -256 350 -252
rect 269 -281 273 -277
rect 306 -285 310 -281
rect 386 -242 390 -238
rect 378 -256 382 -252
rect 415 -260 419 -256
rect 362 -270 366 -266
rect 370 -277 374 -273
rect 399 -277 403 -273
rect 338 -283 342 -279
rect 253 -295 257 -291
rect 261 -302 265 -298
rect 290 -302 294 -298
rect 229 -308 233 -304
rect 330 -305 334 -301
rect 237 -315 241 -311
rect 229 -326 233 -322
rect 269 -315 273 -311
rect 244 -325 248 -321
rect 346 -290 350 -286
rect 378 -290 382 -286
rect 353 -300 357 -296
rect 259 -326 263 -322
rect 277 -325 281 -321
rect 301 -332 305 -325
rect 368 -301 372 -297
rect 386 -300 390 -296
rect 410 -307 414 -300
<< metal2 >>
rect 229 -304 233 -208
rect 237 -311 241 -281
rect 237 -319 241 -315
rect 245 -298 249 -267
rect 253 -291 257 -208
rect 284 -267 288 -263
rect 245 -301 261 -298
rect 245 -321 249 -301
rect 269 -311 273 -281
rect 269 -319 273 -315
rect 277 -294 281 -267
rect 338 -279 342 -207
rect 301 -285 306 -281
rect 277 -297 294 -294
rect 233 -325 244 -322
rect 248 -325 249 -321
rect 277 -321 281 -297
rect 290 -298 294 -297
rect 263 -325 277 -322
rect 301 -325 305 -285
rect 346 -286 350 -256
rect 346 -294 350 -290
rect 354 -273 358 -242
rect 362 -266 366 -207
rect 393 -242 397 -238
rect 354 -276 370 -273
rect 354 -296 358 -276
rect 378 -286 382 -256
rect 378 -294 382 -290
rect 386 -269 390 -242
rect 415 -261 419 -260
rect 410 -265 419 -261
rect 386 -272 403 -269
rect 330 -300 353 -297
rect 357 -300 358 -296
rect 386 -296 390 -272
rect 399 -273 403 -272
rect 330 -301 334 -300
rect 372 -300 386 -297
rect 410 -300 414 -265
<< labels >>
rlabel metal2 338 -208 342 -207 1 ClkB
rlabel metal2 362 -208 366 -207 1 Clk
rlabel metal1 322 -234 323 -211 1 Vpos
rlabel metal1 424 -234 425 -211 1 Vpos
rlabel metal1 322 -344 324 -317 1 Vneg
rlabel metal1 314 -344 316 -317 1 Vneg
rlabel metal1 423 -344 425 -317 1 Vneg
rlabel pwell 213 -344 215 -317 3 Vneg
rlabel metal1 315 -234 316 -211 1 Vpos
rlabel metal1 213 -234 214 -211 3 Vpos
rlabel metal1 312 -311 313 -288 1 Qb
rlabel metal1 421 -311 422 -288 1 Qb
rlabel metal1 312 -285 313 -262 1 Q
rlabel metal1 421 -285 422 -262 1 Q
rlabel metal2 229 -209 233 -208 1 ClkB
rlabel metal2 253 -209 257 -208 1 Clk
rlabel metal1 242 -209 246 -208 1 RstB
rlabel metal1 355 -344 359 -343 1 RST
rlabel metal1 324 -311 325 -262 1 D
rlabel metal1 215 -308 216 -259 3 D
<< end >>
