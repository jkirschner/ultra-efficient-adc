magic
tech scmos
timestamp 1355458399
<< ntransistor >>
rect 12 -6 15 -1
rect 21 -6 24 -1
rect 33 -6 36 -1
rect 90 -6 93 -1
rect 102 -6 105 -1
rect 111 -6 114 -1
<< ptransistor >>
rect 3 49 6 55
rect 19 49 32 76
rect 38 49 41 55
rect 85 49 88 55
rect 94 49 107 76
rect 120 49 123 55
rect 3 22 6 27
rect 21 22 24 27
rect 33 22 36 27
rect 90 22 93 27
rect 102 22 105 27
rect 120 22 123 27
<< ndiffusion >>
rect 11 -5 12 -1
rect 9 -6 12 -5
rect 15 -5 16 -1
rect 20 -5 21 -1
rect 15 -6 21 -5
rect 24 -2 33 -1
rect 24 -6 28 -2
rect 32 -6 33 -2
rect 36 -5 37 -1
rect 89 -5 90 -1
rect 36 -6 39 -5
rect 87 -6 90 -5
rect 93 -2 102 -1
rect 93 -6 94 -2
rect 98 -6 102 -2
rect 105 -5 106 -1
rect 110 -5 111 -1
rect 105 -6 111 -5
rect 114 -5 115 -1
rect 114 -6 117 -5
<< pdiffusion >>
rect 16 55 19 76
rect 0 53 3 55
rect 2 49 3 53
rect 6 54 19 55
rect 6 50 7 54
rect 16 50 19 54
rect 6 49 19 50
rect 32 55 35 76
rect 91 55 94 76
rect 32 51 33 55
rect 37 51 38 55
rect 32 49 38 51
rect 41 51 42 55
rect 84 51 85 55
rect 41 49 44 51
rect 82 49 85 51
rect 88 51 89 55
rect 93 51 94 55
rect 88 49 94 51
rect 107 55 110 76
rect 107 54 120 55
rect 107 50 110 54
rect 119 50 120 54
rect 107 49 120 50
rect 123 53 126 55
rect 123 49 124 53
rect 0 26 3 27
rect 2 22 3 26
rect 6 26 21 27
rect 6 22 16 26
rect 20 22 21 26
rect 24 26 33 27
rect 24 22 26 26
rect 30 22 33 26
rect 36 26 39 27
rect 87 26 90 27
rect 36 22 37 26
rect 89 22 90 26
rect 93 26 102 27
rect 93 22 96 26
rect 100 22 102 26
rect 105 26 120 27
rect 105 22 106 26
rect 110 22 120 26
rect 123 26 126 27
rect 123 22 124 26
<< ndcontact >>
rect 7 -5 11 -1
rect 16 -5 20 -1
rect 28 -6 32 -2
rect 37 -5 41 -1
rect 85 -5 89 -1
rect 94 -6 98 -2
rect 106 -5 110 -1
rect 115 -5 119 -1
<< pdcontact >>
rect -2 49 2 53
rect 7 50 16 54
rect 33 51 37 55
rect 42 51 46 55
rect 80 51 84 55
rect 89 51 93 55
rect 110 50 119 54
rect 124 49 128 53
rect -2 22 2 26
rect 16 22 20 26
rect 26 22 30 26
rect 37 22 41 26
rect 85 22 89 26
rect 96 22 100 26
rect 106 22 110 26
rect 124 22 128 26
<< polysilicon >>
rect 19 77 20 78
rect 24 77 32 78
rect 19 76 32 77
rect 94 77 102 78
rect 106 77 107 78
rect 94 76 107 77
rect 4 56 6 60
rect 3 55 6 56
rect 38 55 41 57
rect 85 55 88 57
rect 120 56 122 60
rect 120 55 123 56
rect 3 47 6 49
rect 19 47 32 49
rect 38 48 41 49
rect 85 48 88 49
rect 94 47 107 49
rect 120 47 123 49
rect 4 28 6 32
rect 23 29 24 33
rect 3 27 6 28
rect 21 27 24 29
rect 33 27 36 29
rect 90 27 93 29
rect 102 29 103 33
rect 102 27 105 29
rect 120 28 122 32
rect 120 27 123 28
rect 3 20 6 22
rect 21 19 24 22
rect 33 20 36 22
rect 90 20 93 22
rect 102 19 105 22
rect 120 20 123 22
rect 21 15 23 19
rect 103 15 105 19
rect 24 1 36 3
rect 12 -1 15 1
rect 21 0 36 1
rect 21 -1 24 0
rect 33 -1 36 0
rect 90 1 102 3
rect 90 0 105 1
rect 90 -1 93 0
rect 102 -1 105 0
rect 111 -1 114 1
rect 12 -7 15 -6
rect 13 -11 15 -7
rect 21 -8 24 -6
rect 33 -8 36 -6
rect 90 -8 93 -6
rect 102 -8 105 -6
rect 111 -7 114 -6
rect 111 -11 113 -7
<< polycontact >>
rect 20 77 24 81
rect 102 77 106 81
rect 0 56 4 60
rect 122 56 126 60
rect 37 44 41 48
rect 85 44 89 48
rect 0 28 4 32
rect 19 29 23 33
rect 33 29 37 33
rect 89 29 93 33
rect 103 29 107 33
rect 122 28 126 32
rect 23 15 27 19
rect 99 15 103 19
rect 20 1 24 5
rect 102 1 106 5
rect 9 -11 13 -7
rect 113 -11 117 -7
<< metal1 >>
rect -13 88 142 102
rect -13 84 -2 88
rect 2 84 124 88
rect 128 84 142 88
rect -13 77 20 81
rect 24 77 102 81
rect 106 77 142 81
rect -2 60 16 64
rect -2 56 0 60
rect -2 53 2 56
rect 7 54 16 60
rect 33 60 93 64
rect 33 55 37 60
rect 89 55 93 60
rect 46 51 80 55
rect 110 60 128 64
rect 110 54 119 60
rect 126 56 128 60
rect -13 44 -10 48
rect -13 36 -10 40
rect -13 29 -10 33
rect -2 32 2 49
rect 44 41 48 51
rect 26 37 48 41
rect 78 41 82 51
rect 124 53 128 56
rect 78 37 100 41
rect -2 28 0 32
rect -2 26 2 28
rect 26 26 30 37
rect 96 26 100 37
rect 124 32 128 49
rect 126 28 128 32
rect 124 26 128 28
rect 41 22 85 26
rect 16 9 20 22
rect 16 -1 20 5
rect 37 -1 41 22
rect 85 12 89 22
rect 121 14 142 18
rect 121 12 129 14
rect 54 5 72 9
rect 85 8 129 12
rect 7 -7 11 -5
rect 85 -1 89 8
rect 137 5 142 9
rect 106 -1 110 1
rect 7 -8 9 -7
rect -13 -11 9 -8
rect 28 -8 32 -6
rect 94 -8 98 -6
rect 115 -7 119 -5
rect 13 -11 113 -8
rect 117 -8 119 -7
rect 117 -11 142 -8
rect -13 -34 142 -11
<< m2contact >>
rect -2 84 2 88
rect 124 84 128 88
rect -2 64 2 68
rect 124 64 128 68
rect -10 44 -6 48
rect -10 36 -6 40
rect -10 29 -6 33
rect 33 44 37 48
rect 89 44 93 48
rect 15 29 19 33
rect 37 29 41 33
rect 85 29 89 33
rect 107 29 111 33
rect 27 15 31 19
rect 16 5 20 9
rect 95 15 99 19
rect 106 18 110 22
rect 50 5 54 9
rect 72 5 76 9
rect 133 5 137 9
rect 106 1 110 5
<< metal2 >>
rect -2 68 2 84
rect 124 68 128 84
rect -6 44 33 48
rect 37 44 89 48
rect 93 44 136 48
rect -6 36 41 40
rect 33 33 41 36
rect 85 36 136 40
rect 85 33 93 36
rect -6 29 15 33
rect 41 29 85 33
rect 111 29 139 33
rect 31 15 95 19
rect 106 9 110 18
rect 20 5 50 9
rect 76 5 133 9
<< labels >>
rlabel metal1 133 16 133 16 1 V+
rlabel metal2 132 6 132 6 1 V-
rlabel metal1 16 -15 16 -15 1 Gnd
rlabel metal1 10 88 10 88 5 Vdd
rlabel metal1 -7 79 -7 79 4 Bias
rlabel m2contact -8 46 -8 46 3 Cascode
rlabel m2contact -8 39 -8 39 3 Thresh
rlabel metal1 -12 30 -12 30 3 Input
<< end >>
