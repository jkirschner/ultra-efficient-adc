* SPICE3 file created from doubleBiasGen.ext - technology: scmos


* Top level circuit doubleBiasGen

M1000 a_38_n9# PosA PosA PosA pfet w=8.1u l=3.9u
+ ad=29.16p pd=39.6u as=68.58p ps=154.8u 
M1001 PosA Bias a_38_n9# PosA pfet w=8.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1002 a_146_n9# Bias PosA PosA pfet w=8.1u l=3.9u
+ ad=29.16p pd=39.6u as=0p ps=0u 
M1003 PosA PosA a_146_n9# PosA pfet w=8.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1004 Cascode PosA PosA PosA pfet w=8.1u l=3.9u
+ ad=29.16p pd=39.6u as=0p ps=0u 
M1005 a_38_n9# Cascode Cascode PosA pfet w=8.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1006 Bias Bias a_38_n9# PosA pfet w=8.1u l=0.9u
+ ad=16.02p pd=38.4u as=0p ps=0u 
M1007 PosA Bias a_1_n53# PosA pfet w=1.8u l=3.9u
+ ad=0p pd=0u as=4.68p ps=13.2u 
M1008 a_79_n61# Bias PosA PosA pfet w=8.1u l=3.9u
+ ad=14.58p pd=19.8u as=0p ps=0u 
M1009 PosA Bias a_79_n61# PosA pfet w=8.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1010 a_1_n53# Bias PosA PosA pfet w=1.8u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1011 a_146_n9# Bias Bias PosA pfet w=8.1u l=0.9u
+ ad=0p pd=0u as=0p ps=0u 
M1012 Cascode Cascode a_146_n9# PosA pfet w=8.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1013 PosA PosA Cascode PosA pfet w=8.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1014 Cascode Vneg Vneg Vneg nfet w=2.1u l=3.9u
+ ad=7.56p pd=15.6u as=16.2p ps=44.4u 
M1015 Vneg a_1_n53# Cascode Vneg nfet w=2.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1016 Bias a_1_n53# Vneg Vneg nfet w=0.9u l=8.1u
+ ad=3.42p pd=10.8u as=0p ps=0u 
M1017 a_73_n59# a_1_n53# a_1_n53# Vneg nfet w=8.1u l=3.9u
+ ad=11.79p pd=27u as=16.02p ps=38.4u 
M1018 a_1_n53# a_1_n53# a_111_n59# Vneg nfet w=8.1u l=3.9u
+ ad=0p pd=0u as=11.79p ps=27u 
M1019 Vneg a_1_n53# Bias Vneg nfet w=0.9u l=8.1u
+ ad=0p pd=0u as=0p ps=0u 
M1020 Cascode a_1_n53# Vneg Vneg nfet w=2.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1021 Vneg Vneg Cascode Vneg nfet w=2.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1022 a_73_n59# a_1_n53# Vneg Vneg nfet w=2.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1023 a_79_n61# a_79_n61# a_73_n59# Vneg nfet w=2.1u l=3.9u
+ ad=3.78p pd=7.8u as=0p ps=0u 
M1024 a_111_n59# a_79_n61# a_79_n61# Vneg nfet w=2.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
M1025 Vneg a_1_n53# a_111_n59# Vneg nfet w=2.1u l=3.9u
+ ad=0p pd=0u as=0p ps=0u 
C0 Vneg gnd! 6.4fFCascodeC1 PosA gnd! 7.5fFCascodeC2 a_79_n61# gnd! 4.5fFVnegC3 a_1_n53# gnd! 2.0fFCascodeC4 Vneg gnd! 3.5fFBiasC5 PosA gnd! 23.0fFBiasC6 a_1_n53# gnd! 12.3fFVnegC7 a_1_n53# gnd! 2.3fFPosA.end

