magic
tech scmos
timestamp 1355754911
<< error_s >>
rect 361 3997 372 4000
rect 361 3996 400 3997
rect 361 3523 372 3526
rect 361 3522 400 3523
rect 361 3049 372 3052
rect 361 3048 400 3049
rect 507 2979 513 2980
rect 4636 2734 4998 2735
rect 361 1153 372 1156
rect 361 1152 400 1153
<< metal1 >>
rect 575 4481 579 4487
rect 596 4481 599 4487
rect 575 4476 599 4481
rect 602 4465 606 4488
rect 1049 4481 1053 4487
rect 1070 4481 1073 4487
rect 1049 4476 1073 4481
rect 1076 4471 1080 4488
rect 1523 4481 1527 4491
rect 1544 4481 1547 4490
rect 1523 4476 1547 4481
rect 510 4394 554 4398
rect 513 4388 526 4391
rect 521 4371 526 4388
rect 513 4367 526 4371
rect 541 4022 554 4394
rect 596 4105 609 4465
rect 1033 4464 1080 4471
rect 1550 4464 1554 4487
rect 596 4080 986 4105
rect 541 3997 935 4022
rect 541 3924 879 3945
rect 509 3920 879 3924
rect 513 3914 526 3917
rect 521 3897 526 3914
rect 513 3893 526 3897
rect 551 3450 840 3461
rect 509 3446 840 3450
rect 513 3440 526 3443
rect 521 3423 526 3440
rect 513 3419 526 3423
rect 828 3267 840 3446
rect 860 3416 879 3920
rect 914 3563 935 3997
rect 969 3717 986 4080
rect 1033 3868 1050 4464
rect 1550 4447 1701 4464
rect 1681 4016 1701 4447
rect 1921 4139 1947 4494
rect 2018 4186 2034 4492
rect 2479 4417 2488 4491
rect 2437 4400 2488 4417
rect 2018 4160 2322 4186
rect 2307 4135 2322 4160
rect 2437 4151 2472 4400
rect 2493 4162 2508 4491
rect 2945 4483 2949 4487
rect 2966 4483 2969 4487
rect 2945 4479 2969 4483
rect 2972 4456 2976 4489
rect 3419 4482 3423 4487
rect 3440 4482 3443 4487
rect 3419 4477 3443 4482
rect 3446 4476 3450 4492
rect 3572 4482 3579 4485
rect 3582 4482 3591 4485
rect 2972 4452 2973 4456
rect 3446 4387 3454 4476
rect 3568 4473 3571 4476
rect 3574 4473 3577 4482
rect 3568 4470 3577 4473
rect 3582 4479 3585 4482
rect 3588 4479 3591 4482
rect 3582 4476 3591 4479
rect 3582 4470 3585 4476
rect 3588 4470 3591 4476
rect 3594 4482 3604 4485
rect 3594 4479 3597 4482
rect 3600 4479 3604 4482
rect 3607 4482 3613 4485
rect 3616 4484 3625 4485
rect 3616 4482 3626 4484
rect 3607 4479 3610 4482
rect 3594 4476 3603 4479
rect 3607 4476 3613 4479
rect 3594 4470 3597 4476
rect 3600 4470 3604 4476
rect 3607 4473 3610 4476
rect 3616 4473 3619 4482
rect 3622 4481 3626 4482
rect 3623 4474 3626 4481
rect 3640 4482 3650 4485
rect 3653 4482 3662 4485
rect 3640 4479 3643 4482
rect 3653 4479 3656 4482
rect 3659 4479 3662 4482
rect 3640 4476 3650 4479
rect 3622 4473 3626 4474
rect 3646 4473 3650 4476
rect 3607 4470 3613 4473
rect 3616 4471 3626 4473
rect 3616 4470 3625 4471
rect 3630 4470 3634 4473
rect 3640 4470 3650 4473
rect 3653 4476 3662 4479
rect 3653 4470 3656 4476
rect 3659 4470 3662 4476
rect 3665 4482 3682 4485
rect 3665 4470 3668 4482
rect 3672 4470 3675 4482
rect 3679 4470 3682 4482
rect 3693 4482 3702 4485
rect 3693 4479 3696 4482
rect 3699 4479 3702 4482
rect 3693 4476 3702 4479
rect 3686 4470 3690 4473
rect 3693 4470 3696 4476
rect 3699 4470 3702 4476
rect 3705 4482 3722 4485
rect 3705 4470 3708 4482
rect 3712 4470 3715 4482
rect 3719 4470 3722 4482
rect 3725 4479 3728 4485
rect 3731 4479 3734 4485
rect 3725 4476 3734 4479
rect 3728 4470 3731 4476
rect 3631 4468 3634 4470
rect 3687 4468 3690 4470
rect 4464 4394 4491 4398
rect 2492 4140 2561 4162
rect 1681 3999 1684 4016
rect 1700 3999 1701 4016
rect 4479 3947 4487 3951
rect 4479 3930 4483 3947
rect 4479 3927 4487 3930
rect 1033 3866 1700 3868
rect 1033 3851 1684 3866
rect 969 3700 1688 3717
rect 1700 3700 1702 3717
rect 914 3548 1688 3563
rect 4479 3473 4487 3477
rect 4479 3456 4483 3473
rect 4479 3453 4487 3456
rect 4468 3447 4488 3450
rect 4472 3446 4488 3447
rect 4472 3443 4475 3446
rect 860 3401 1687 3416
rect 861 3400 1702 3401
rect 828 3251 1688 3267
rect 1470 3101 1683 3117
rect 1697 3101 1698 3117
rect 1470 2987 1485 3101
rect 552 2977 1485 2987
rect 510 2972 1485 2977
rect 513 2966 526 2969
rect 1506 2967 1698 2968
rect 521 2949 526 2966
rect 513 2945 526 2949
rect 1505 2952 1682 2967
rect 1697 2952 1698 2967
rect 4339 2966 4492 2982
rect 1505 2513 1524 2952
rect 547 2502 1524 2513
rect 509 2498 1524 2502
rect 1559 2805 1683 2820
rect 513 2492 526 2495
rect 521 2475 526 2492
rect 513 2471 526 2475
rect 1559 2040 1580 2805
rect 1513 2039 1580 2040
rect 547 2028 1580 2039
rect 511 2024 1580 2028
rect 1615 2654 1685 2671
rect 1697 2654 1698 2671
rect 513 2018 526 2021
rect 521 2001 526 2018
rect 513 1997 526 2001
rect 1615 1565 1638 2654
rect 4339 2375 4370 2966
rect 3480 2349 4370 2375
rect 4389 2493 4491 2509
rect 3480 2348 4365 2349
rect 4389 2338 4417 2493
rect 3479 2310 4417 2338
rect 3137 1976 3614 1981
rect 3137 1922 3141 1976
rect 531 1554 1638 1565
rect 510 1550 1638 1554
rect 1615 1549 1638 1550
rect 510 1544 526 1547
rect 521 1527 526 1544
rect 509 1523 526 1527
rect 508 1076 570 1080
rect 509 1070 529 1073
rect 525 1053 529 1070
rect 509 1049 529 1053
rect 564 1060 570 1076
rect 564 1045 1664 1060
rect 562 906 1664 921
rect 562 611 588 906
rect 1056 905 1664 906
rect 1803 796 1836 880
rect 520 606 588 611
rect 509 602 588 606
rect 700 770 1836 796
rect 512 596 525 599
rect 521 579 525 596
rect 509 575 525 579
rect 700 544 726 770
rect 2386 715 2400 857
rect 596 528 726 544
rect 1534 689 2400 715
rect 596 512 612 528
rect 1534 526 1560 689
rect 3588 611 3614 1976
rect 4480 1103 4487 1107
rect 4480 1086 4483 1103
rect 4480 1083 4487 1086
rect 4446 1076 4488 1080
rect 4446 1066 4472 1076
rect 4480 629 4491 633
rect 4480 612 4483 629
rect 3588 606 4472 611
rect 4480 609 4487 612
rect 3588 602 4493 606
rect 3588 598 4472 602
rect 3588 585 4446 598
rect 1550 513 1554 526
rect 1557 516 1581 520
rect 1557 513 1560 516
rect 1577 513 1581 516
rect 2031 516 2055 519
rect 2031 513 2034 516
rect 2051 513 2055 516
rect 2505 516 2529 519
rect 2505 513 2508 516
rect 2525 513 2529 516
rect 2979 516 3003 519
rect 2979 513 2982 516
rect 2999 513 3003 516
rect 3453 516 3477 519
rect 3453 513 3456 516
rect 3473 513 3477 516
rect 3927 516 3951 519
rect 3927 513 3930 516
rect 3947 513 3951 516
rect 4394 511 4398 516
rect 4401 516 4425 519
rect 4401 511 4404 516
rect 4421 513 4425 516
<< m2contact >>
rect 2973 4452 2979 4456
rect 3446 4373 3454 4387
rect 1684 3999 1700 4016
rect 4487 3920 4492 3924
rect 1684 3850 1700 3866
rect 1688 3700 1700 3717
rect 1688 3548 1702 3563
rect 4468 3443 4472 3447
rect 1687 3401 1702 3416
rect 1688 3251 1702 3267
rect 1683 3101 1697 3117
rect 1682 2952 1697 2967
rect 1683 2805 1697 2820
rect 1685 2654 1697 2671
rect 2389 2077 2393 2082
rect 2988 1885 2992 1889
rect 1664 1045 1674 1060
rect 1664 905 1674 921
rect 3433 853 3455 859
rect 4433 1066 4446 1080
rect 2024 513 2028 517
rect 2498 513 2502 517
rect 2972 513 2976 517
rect 3446 513 3450 517
rect 3920 513 3924 517
rect 4394 516 4398 520
<< metal2 >>
rect 2973 4450 2979 4452
rect 2973 4435 2974 4450
rect 2978 4435 2979 4450
rect 2973 4434 2979 4435
rect 4481 3920 4487 3924
rect 1687 3563 1702 3564
rect 1687 3548 1688 3563
rect 4467 3443 4468 3447
rect 1687 3400 1702 3401
rect 4451 2018 4452 2034
rect 4456 2018 4491 2034
rect 4451 2017 4491 2018
rect 3198 1954 3202 1956
rect 3198 1948 3549 1954
rect 3198 1937 3202 1948
rect 3523 1079 3549 1948
rect 4484 1545 4489 1559
rect 3523 1053 4433 1079
rect 2608 754 2633 859
rect 1070 728 2633 754
rect 1070 509 1086 728
<< m3contact >>
rect 2974 4435 2978 4450
rect 3446 4359 3454 4373
rect 4477 3920 4481 3924
rect 4463 3443 4467 3447
rect 2389 2072 2393 2077
rect 4452 2018 4456 2034
rect 3079 1885 3083 1889
rect 2379 1706 2394 1718
rect 4480 1545 4484 1559
rect 3433 847 3455 853
rect 2024 517 2028 521
rect 2498 517 2502 521
rect 2972 517 2976 521
rect 3446 517 3450 521
rect 3920 517 3924 521
rect 4394 520 4398 524
<< metal3 >>
rect 2586 4450 2979 4452
rect 2586 4435 2974 4450
rect 2978 4435 2979 4450
rect 2586 4434 2979 4435
rect 2586 2411 2603 4434
rect 2620 4373 3456 4376
rect 2620 4359 3446 4373
rect 3454 4359 3456 4373
rect 2620 4357 3456 4359
rect 2620 2501 2637 4357
rect 3558 3924 4483 3926
rect 3558 3920 4477 3924
rect 4481 3920 4483 3924
rect 3558 3918 4483 3920
rect 3558 3901 4473 3918
rect 2620 2488 2638 2501
rect 2590 2078 2601 2411
rect 2388 2077 2601 2078
rect 2388 2072 2389 2077
rect 2393 2072 2601 2077
rect 2388 2071 2600 2072
rect 2621 1720 2638 2488
rect 3558 1912 3584 3901
rect 2983 1904 3584 1912
rect 3652 3447 4470 3450
rect 3652 3443 4463 3447
rect 4467 3443 4470 3447
rect 3652 3425 4470 3443
rect 2983 1903 3574 1904
rect 2983 1885 2990 1903
rect 3652 1892 3678 3425
rect 3077 1889 3678 1892
rect 3077 1885 3079 1889
rect 3083 1885 3678 1889
rect 2983 1884 2989 1885
rect 3077 1883 3678 1885
rect 3900 2034 4459 2041
rect 3900 2018 4452 2034
rect 4456 2018 4459 2034
rect 3900 2015 4459 2018
rect 3900 1833 3926 2015
rect 3497 1807 3926 1833
rect 3497 1768 3926 1794
rect 2378 1718 2638 1720
rect 2378 1706 2379 1718
rect 2394 1706 2638 1718
rect 2378 1705 2638 1706
rect 2379 1704 2638 1705
rect 3900 1560 3926 1768
rect 3900 1559 4487 1560
rect 3900 1545 4480 1559
rect 4484 1545 4487 1559
rect 4452 1544 4487 1545
rect 649 864 682 865
rect 649 829 1784 864
rect 649 799 682 829
rect 648 750 682 799
rect 2522 793 2548 897
rect 2015 767 2548 793
rect 648 571 681 750
rect 520 570 681 571
rect 519 551 681 570
rect 519 532 532 551
rect 491 493 532 532
rect 2015 521 2041 767
rect 2639 702 2665 897
rect 2015 520 2024 521
rect 2023 517 2024 520
rect 2028 520 2041 521
rect 2483 676 2665 702
rect 2756 702 2782 897
rect 2938 741 2964 897
rect 3042 780 3068 897
rect 3198 819 3224 897
rect 3432 853 3456 854
rect 3432 847 3433 853
rect 3455 847 3588 853
rect 3432 846 3588 847
rect 3433 833 3588 846
rect 3614 833 4462 853
rect 3198 793 3588 819
rect 3614 793 4407 819
rect 3042 754 3588 780
rect 3614 754 3926 780
rect 2938 715 3458 741
rect 2756 676 2977 702
rect 2483 521 2509 676
rect 2483 520 2498 521
rect 2028 517 2029 520
rect 2023 516 2029 517
rect 2497 517 2498 520
rect 2502 520 2509 521
rect 2951 521 2977 676
rect 2951 520 2972 521
rect 2502 517 2503 520
rect 2497 516 2503 517
rect 2971 517 2972 520
rect 2976 517 2977 521
rect 3432 521 3458 715
rect 3432 520 3446 521
rect 2971 516 2977 517
rect 3445 517 3446 520
rect 3450 520 3458 521
rect 3900 521 3926 754
rect 3900 520 3920 521
rect 3450 517 3451 520
rect 3445 516 3451 517
rect 3919 517 3920 520
rect 3924 520 3926 521
rect 4381 524 4407 793
rect 4381 520 4394 524
rect 4398 520 4407 524
rect 4439 533 4461 833
rect 3924 517 3925 520
rect 4387 519 4399 520
rect 4439 519 4528 533
rect 3919 516 3925 517
rect 4515 407 4528 519
rect 4593 414 4594 419
rect 4518 401 4528 407
use iopad  iopad_10
timestamp 1259953556
transform -1 0 841 0 -1 5000
box -2 0 476 513
use iopad  iopad_11
timestamp 1259953556
transform -1 0 1315 0 -1 5000
box -2 0 476 513
use iopad  iopad_12
timestamp 1259953556
transform -1 0 1789 0 -1 5000
box -2 0 476 513
use inpad  inpad_2
timestamp 1259953556
transform -1 0 2263 0 -1 5000
box -2 0 476 513
use inpad  inpad_3
timestamp 1259953556
transform -1 0 2737 0 -1 5000
box -2 0 476 513
use iopad  iopad_22
timestamp 1259953556
transform -1 0 3211 0 -1 5000
box -2 0 476 513
use iopad  iopad_23
timestamp 1259953556
transform -1 0 3685 0 -1 5000
box -2 0 476 513
use blankpad  blankpad_10
timestamp 1259953556
transform -1 0 4159 0 -1 5000
box -2 0 476 513
use blankpad  blankpad_9
timestamp 1259953556
transform -1 0 4633 0 -1 5000
box -2 0 476 513
use padframe_top  padframe_top_0
timestamp 1259953556
transform 1 0 0 0 1 4487
box 0 0 5000 513
use iopad  iopad_1
timestamp 1259953556
transform 0 1 0 -1 0 4633
box -2 0 476 513
use iopad  iopad_0
timestamp 1259953556
transform 0 -1 5000 1 0 4159
box -2 0 476 513
use iopad  iopad_2
timestamp 1259953556
transform 0 1 0 -1 0 4159
box -2 0 476 513
use iopad  iopad_3
timestamp 1259953556
transform 0 1 0 -1 0 3685
box -2 0 476 513
use iopad  iopad_4
timestamp 1259953556
transform 0 1 0 -1 0 3211
box -2 0 476 513
use iopad  iopad_5
timestamp 1259953556
transform 0 1 0 -1 0 2737
box -2 0 476 513
use iopad  iopad_6
timestamp 1259953556
transform 0 1 0 -1 0 2263
box -2 0 476 513
use iopad  iopad_7
timestamp 1259953556
transform 0 1 0 -1 0 1789
box -2 0 476 513
use OverallLayout_FINAL  OverallLayout_FINAL_0
timestamp 1355723001
transform -1 0 2182 0 -1 4069
box -1328 -86 518 3217
use iopad  iopad_25
timestamp 1259953556
transform 0 -1 5000 1 0 3685
box -2 0 476 513
use iopad  iopad_24
timestamp 1259953556
transform 0 -1 5000 1 0 3211
box -2 0 476 513
use inorpad  inorpad_3
timestamp 1259953556
transform 0 -1 5000 1 0 2737
box -2 0 476 513
use inorpad  inorpad_2
timestamp 1259953556
transform 0 -1 5000 1 0 2264
box -2 0 476 513
use inorpad  inorpad_1
timestamp 1259953556
transform 0 -1 5000 1 0 1789
box -2 0 476 513
use inorpad  inorpad_0
timestamp 1259953556
transform 0 -1 5000 1 0 1315
box -2 0 476 513
use iopad  iopad_8
timestamp 1259953556
transform 0 1 0 -1 0 1315
box -2 0 476 513
use iopad  iopad_21
timestamp 1259953556
transform 0 -1 5000 1 0 841
box -2 0 476 513
use padframe_left  padframe_left_0
timestamp 1259953556
transform 1 0 0 0 1 367
box 2 2 513 4264
use iopad  iopad_9
timestamp 1259953556
transform 0 1 0 -1 0 841
box -2 0 476 513
use inpad  inpad_0
timestamp 1259953556
transform 1 0 367 0 1 0
box -2 0 476 513
use inpad  inpad_1
timestamp 1259953556
transform 1 0 841 0 1 0
box -2 0 476 513
use iopad  iopad_19
timestamp 1259953556
transform 1 0 1315 0 1 0
box -2 0 476 513
use iopad  iopad_18
timestamp 1259953556
transform 1 0 1789 0 1 0
box -2 0 476 513
use iopad  iopad_17
timestamp 1259953556
transform 1 0 2263 0 1 0
box -2 0 476 513
use iopad  iopad_16
timestamp 1259953556
transform 1 0 2737 0 1 0
box -2 0 476 513
use iopad  iopad_15
timestamp 1259953556
transform 1 0 3211 0 1 0
box -2 0 476 513
use iopad  iopad_14
timestamp 1259953556
transform 1 0 3685 0 1 0
box -2 0 476 513
use padframe_right  padframe_right_0
timestamp 1259953556
transform 1 0 4487 0 1 367
box 0 2 511 4264
use iopad  iopad_20
timestamp 1259953556
transform 0 -1 5000 1 0 367
box -2 0 476 513
use iopad  iopad_13
timestamp 1259953556
transform 1 0 4159 0 1 0
box -2 0 476 513
use padframe_bottom  padframe_bottom_0
timestamp 1259953556
transform 1 0 0 0 1 0
box 0 0 5000 513
<< labels >>
rlabel m2contact 1701 3258 1701 3258 1 Bit8
rlabel m2contact 1699 3407 1699 3407 1 Bit9
rlabel m2contact 1697 3555 1697 3555 1 Bit10
rlabel space 1061 4487 1061 4487 8 Bias
rlabel space 587 4487 587 4487 8 Bias
rlabel space 4487 1094 4487 1094 4 Bias
rlabel metal2 4387 1069 4387 1069 1 CLC2
rlabel metal1 4354 594 4354 594 1 CLC1
rlabel metal3 4444 2028 4444 2028 1 Iref
rlabel space 4487 3938 4487 3938 4 Bias
rlabel metal3 3672 1909 3672 1909 1 Shunt_Iin
rlabel metal3 3571 2019 3571 2019 1 Shunt_Iref
<< end >>
